library ieee;
use ieee.std_logic_1164.all;


entity lfsr_13bit is

end entity lfsr_13bit;


architecture behaviour of lfsr_13bit is

begin

end architecture behaviour;

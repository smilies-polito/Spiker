library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rf_signed_tb is
end entity rf_signed_tb;

architecture test of rf_signed_tb is

begin

end architecture test;

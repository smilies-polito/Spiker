library ieee;
use ieee.std_logic_1164.all;

entity spiker is

end entity spiker;

architecture behaviour of spiker is

begin


end architecture behaviour;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity shifter is

	port(
				
	);

end entity shifter;


architecture behaviour of shifter is
begin

end architecture behaviour;

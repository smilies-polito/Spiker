library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity layer_datapath is

end entoty layer_datapath;


architecture behaviour of layer_datapath is

begin


end architecture behaviour;

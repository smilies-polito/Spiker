library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_784x128_exc_ip is
	port(
		clka	: in std_logic;
		addra	: in std_logic_vector(9 downto 0);
		douta	: out std_logic_vector(511 downto 0)
	);
end entity rom_784x128_exc_ip; 

architecture behavior of rom_784x128_exc_ip is

	type rom_type is array(0 to 783) of std_logic_vector(511 downto 0);

	constant mem	: rom_type := (
		
		"01110111011101110111000001110000011100110111000001000011011101100111011100010011000101110101010001000010001000100011000001110000011101110111011101000111000000100111010101110111011100000010011100000111011100110110011101100111011101110101010101110111011101010011011101110110001001110111010000010100011101110111011101110111001000010001011101100111011101110000010000010111001000000111010100000110011100010111011101110100011001000101010101110111011101110101010000010101011101000111000001110100010001100111011101110101",
		"01000011011100010101011100000000011101110100011101110101001101110101011101010000011101110001000000100100011100010000010101000000011101110101000000110111011100100111011100100111011100010110011101110001010101110100011101110010000001010111011101000111001101110001011101110111011101100011011100100111001101110011011101010000011100110100011101110111010001110111001001110111011101110111011101110111000000010000000101110001011101100011011100010111011001110111011001110001011101110111011101110100010001100111011101000111",
		"01110111011101110110010001110101011101110111011101110110000101110111010101110111011100010001011101110010011101110011000001110110011101110110000100100111000001000101011101110110011100000101000001110110011101110111011101110110011101000111011101110111010000010101011101110111011101110101011001100111000000010111011100010111001101100111001101110111011100110101011101110111010101110111001100010011001101110001000101000111010001110111011101110010011101110101000101110101010100110011011101110111011101110111011101000000",
		"00100111011001110010011101000101011101010101011100000000001001000111011101110111000101100111001101110111001000100110001100110111001101100111010001110111011101110111011101110111000100100011010000110111010100010001011001110111001101110110011100010010000101110101001001110100011100010111001001110100000001110000011100000111000001110111010101110111011101100110011101110011010101000010011101100111001001110111011101110110011101110111010001100111000101110110010001110111011101110101011101000111011101010111000001110111",
		"01000111011000010111011101110111011101100111001100010101011101110111011101110010011101100111011101110111011101110111011100110100011101010111011101110000010000000111011101110111001001110111011101110000001101110111000101110111011101110111011100110011011101110111011100110111011101110101011001010111011101110100011100100111011101110011011101000001011101010010010000000111011101110111011101100011011101110001011100000010011100000111011101110001011101100111011101110111010001110111001100010111011000110110011101110010",
		"01110101011101110111010001110111010001110110011101110111011101000011001001110111010100000111011001110111011101110111011100000100011101110111011001010111000101110001001001100010010001110111010001110111011100110111011100100001011101110110011001110101011100000111011101110111011101110110010100100011011101110111010101010110011101110000000101110010000101110101011100100001011101110010001101100111011100110111011101000111000101110000001101100000011001110110011101110101000001110111001101110110011101110111011001010111",
		"01110111011101110111011101110111011101010001011101110111011101010111011101110111011101110100000101110111011101000001011101110000011101110111011101010111001101010111001001110111001101110011011000110011011101110111000101010101011100110010011100100001011101110111011101110011000101110111011100100110011101110111011101110011000001110111011101110000001001110110011101100101010001110111010001110111000000100111011101110111011101110111011100100000010101110111011100010111011101110111011101100111001001110111011101110110",
		"01110111011100000100001000000111011101110111011101100111010101110111011101110111011100100100011101110001001001110000011101110111011101100001001001110111001001110010011101110111001001100111001001110101011101110111011101110110001100010101011100000110011101110010010001110111011100010010011100100010011100000111011101110010011000110111001101110111011000110101011101110100011100010001001101110111010100110111001001000111011101110111011101110011011100000111011101000111011100010111011101110100011001110111011101000101",
		"00100010011100000111011100100100000001110010000101110101011100100111011101110001011101110000001100110111011101110111010101110111011101110111011101110100000101100010011101110100011101110100010001110000011001110111001101110111011101110111011101110100011101010000010101100100011101110111001001110000001000110011011101110111011100000111011101110000011101110111011101110111011101110111011101010011011101010011011101110001001101110111011101110111010101110111001101110001011101110111001001110111011001110110011100000111",
		"00000111011101110111011000100111011100110111000001110111011101110101001101010111011101010111011101110110011101010111011101110010001101110111000101000111011101010111011101110111011100110111010100010000011001110110011101100111011100010000011101000111011101110100001101110111011000000111010000110010011101110111011101110101001100010101011100110111011101000111011101100111011101110110000101110111011101110101011001110010011101110000001001110111011101110110010101110101011101100111011001110111000101110111011101110111",
		"01110011010100100011011100100010011100010110011101110100001001110111001001110110011001110111000101110010010000110111010100100111001101110111011100110011011101110000011101110111011101110111011101110111011000000010011101000111001100100001011101110111001101110111011101110110011101110000011101110111011101110011000001110101001100000111011101110111011101110111011101110000000001110111010101110001011101100011011101110111011101000000001001110101011101100111011101100001011101100011001101110001000101110111000001110111",
		"01110111011101110000011100000010000101010111000101010111011100100111011101110101011100110000011101110111011000110001011101110111010101000010010101110101011101110010010000110111001101110000011001110001011101110000011101110101001000010001011101010111011101010010011100000010011101110110011100100100001100010001011101110111011101110101010100010000011100010111011101110011000100110001011101110111000000100111011001100111011101110011000100010111011100100001011101110001001001110100011101010111011101110111011101110111",
		"00000111011101110111011101010111001101110110011100110111011101010110000101110111011101010000011101110111011100000100000100100101011101000111010001110101011100100111000001110111011100000111010001110000001101100001001101110100011101110111000001000111011101110111011101110111010101110111011101110111011101110111011001110111011101110100011101110010011100010111011101010111011101000111000001010111001001110111011101110111000001110000001101110111011100100110011101100111011101110000011101110001000001110111011101100111",
		"01110111011100010111011101110111011100100111010101010111011100100111011101000011011001110111011100100111011101110111011100000111000000010000010101000111011101110111011100000111010101110010011101000111011100110111001100010111011100000111011101110010011101110100011100100111000101110100011101110111000100010111011101110110000001110001010001000111000001110111011100110111011101110111000001110111011101110111011101110011001001000111011101110111000001110111011101110111000001110101011101110111011100110111011101110010",
		"01110100011101100110011101000100001101100111011101110010011100010111011001110111010000010110011101110111011101100111010101110111011101110000011101110111011101110111010100110111011100000111011101110101011101000111011101110111011101110111010001110111011100110000011101000010001001110111010101100111000101110001011101000111010001010111011101110111010101110110000001110111000101110100010001100010001001000111000101110111011101110110011101000111011100000111011101110100011100000001011101100111001001110111000101100111",
		"00000011011101100111011101010001000101110111011101110110011101110010010101000000011101110110011101110111011100000011001100110111011101110111010101110111011101110011011101110101011101100010001001100111011101110111000100010110010001010100011101110001001001110101001101110000011101110111011101110111011100110110011101010111000001110110011100000101011101110111011101000111011101110111010001010111000000110100011101010111000001110111010000110111011001110111011100100111011101110101000000110000010001000011011101110111",
		"01010111011101010010011101110111000001110101011101110111010000100111010001100010011101110101010000000111011101110111001101110000011101110101001001100111000001110111011101110111011101110111011101110111011101110000001001110111011100010110011101110111011101110111011101110110001001110010011001100111000001110111011001100111010101100111010001110111010101110111011101110111010101110111011100100001000101110111001100100111011101110001000001110100011101100111010101110111011101110010010001100111011101110000011101110000",
		"01110110011101100010001001110111010101110111011101110111011101110100011101110111000101110111011100000011010001110111011101110101001101110000001000000111011101110111011101000111011101110111011101110010011100000110010001110010001101110001001101110111010001110010001101010101011100010111010001110100000000000011011101110111011101110010010101100000011101110111000000100011010101110111001001000000000101000111000101110111011101000111011100100101000001110101011101110100000001110111011101110000000101000111011101110011",
		"00010010011101110111000000110101011101110111011101110000011101110010011100010111011101110111011101110111011101100000001101000101011101110100001100010111011101110000001100000000011100010101011101110111011100010101011000110111010101110000011101110111000000110111011101110111011100110111011101110111000001110111011101110001011101110011011100100111010101110111001101110111011101110111000101110000011101110101011001110001010000010111000101110111011101110111001100010000010000000001010101100001011101110100000101110111",
		"00010111001000110111000101110000011101000111011101110111011101100100011101110111011001100000011100100000011101110000010101110110000101110101011100110111011101100010011100000001000001110111011101110111010101110001011100000011000101110111011101110111011101010111010101110001011101010111011101000000010101000011000101010111011101000011011100110011000001110111011101110011011101110001011101110111011100000111001101110101010101110011011100000010001001110100011101110001000101110111011101110010011100100111011101110111",
		"01010101011101000111011101000111011101010111011101110010010101110111011101110011011101110110011001110111011101110111001101110111011101110101011101110111011101110111010101100111011101110111011101110010011101000111011101110111001000110100011100000011011101100111011101110000011101110111011101010111010001110101011101110000011101110111011101110111011101110111011101110111010101110000011100110111011001110000011101110111011101110111000100000111011101000111010101110100001101110111000001110111011101010100011101110111",
		"01110101011101110111011101110111011100100111011101110111011101000111011101110100011001110011011101100001001101110011000101110000011001000111011101110111011100010100011001110110011000100111011101100101011001110110011100010001010000100110011100100001010001110101011101110101010101000101011100110111011100100011011001010110001000110111011101010111011101110001011101110111011101110111011101110111011101110111010000010000011101110000000100010111011100000000001101110111011101110001011101110001011101110100011101110010",
		"00100111011101110111011101110111011101000111001100100111011100110111011100010000010001110111010001110111001001110110010001110111011101110110011100100111000101110010000100010110011001110101011101110111011100110111011101010001011100110111000101110111011100100111011100000000001100100011001000100100011101110111011101110110000001110111000001100111011001000111000101110010011101110111011101110001011101110101011101110111011001110000011101110111011101110111011101110111011101010111011101110000000100100100010101110111",
		"01110010011101110110000001110011010001110111000000010111001000110111011001110111011101110111011101110111010101100111011101110111010000010111010001110110011101100111011101110111011101110111001101100111010101110111000000000001000101010000001100100100011101110111011101110010001100010110000000110110010101110110011101110101011101110111011101110011011101110011011101110111010001010101010001110111001001010111001101110111000000110111011101110111011101110011001000110111011101110001011101000111010001110111001100010010",
		"00000010011001110001010101000111010001000001011100110111010101000111011101110111011101010011011101110111001001000000010000110010011101110100011101110110011101110111011101110101011100100111011100000111001101110110011101010111010000010111011101010000001001110111010101110100000100010000011101110111011101110111011101110111000001110100011101010110011100100111011101110011011001110111011101110111011101110001011101110111010101110000000001110111011100000001000101110111011101010111010101110111010101110101011101110001",
		"01110111011101110110011101110111011001110111011101100111011100110111011101100111001001110111011001000111011101010111011101110111011101110110011100010111011101110111011101000101000101110010011101110001011100100100011100000011011101010111001100000111011101110101011100010100010100010110011101110010011101010111011001110001010000010001011101110111011100000100010000110111011100100011011100110010011101110111011001110001000101110111011101110111011101110111011100110010001000110111001001110111011101010110000001000110",
		"00100111011101110111000101110111011101110010011101100111011101110111011101000100011101010110011101110001011100110111000101110111000101110111010101110100011101010011011101000111000000000111001101000111010001110111011101000011000101110111001101110111001001110011010101110000011101010001011101110100011100110111011101110000011101100111000001110000001101100110011100000001001101110001011101110111011101100111011100100111011000100100010001110111011101110010011101100111011101110111000100100111011100010111010001100100",
		"00010000011101100111011101010111001001000011011100100111000101100010011101110111011101110111011100110111010001110111010101110011011100100110011101110111011101110011011101110111011100000001011101110010010001110111011101010111001101110111011101110110000100100111001101110111011101110110000101010101001000100111011100110101011100000010011100100101010000000111011101110010011100100110011101110111011100110111010000110001011101110101011101110011001001000011000000100111001001110110000101110111011100110111011100100110",
		"01110111011100110111011101110000011100010110011101110111011101110100011101010100001001000110011100110111001100000001000001110111011101110111011100100111011100110111011101110111011101110111011001110111000100000111011101010111001101110111011101110000011101010111000101100111011101110111011101010111010101110011011101000110011101110111011100100111011001110111010101100011010001110111000100100111011100010110011101000010011101000000011101110110000000100111000001110111011101110111001101110101011101110101011100010100",
		"01110101011101110100000101110011000000110010010000110111011100000011010001110111011101100011010101110111001101110001011001110111011100100100010101100111011101110111010001110011000001110111001000010101011101110101000101110111011101110111011101110111000001110010010101000111011101110111011101000111011101110111011101110010001100010111001101110001010100000110011100000001001100000100001000000000001100010111010100000100011001110111001001110111011101010010011100100111011101110111000001100111001101110100011001110111",
		"01110000011101110101011001110111010001010111011101110101001100110111011101110111011101110000011101010011010101110111011100100111011101110111011001000111011101110000011001110111011101110100000000010000011000100110011101100111011100100100011101110000000001110111011100110111010100100111011101110111010101010100011101110100001101110010011100110111000101110001001001000110011100010000011101110111010101110001001001110111011101110111011100010111011101110000000100000111000000010111001101110111011001000010011101010000",
		"00110000011101100111011101110000001101110111011101110101010000010101011001110111001001110100011100110101001101100111011100100111011101110111001001100111011100100001011001110001011101110000010101110100000001110000011101110100010100110111011101110111011100110111011101110111011101100111001100100000001001110111001001110111011100110100011101110111001100110111011101110111000101110111011101110111011101100111011101110000011101110111011101110100011101110111010000110010001101110111010001010101011100110010011101110011",
		"00100111001001110111001001110111011101110111011101110101000101010011000000110111011101110011010001010111011101000000011101110111000100110000000100100110010001110111011101100111011100010000000001110111011100100111011101110100011101110110010001110111011101110111011101110111001101010111011101010111011101110011010001110110010001110001000100110111011101100000011101110111011101110111011101110001011101000111011101110001011101100010000001110010011101010111011101110111000100000111011101110111001101110111010001110101",
		"01110111011100100111011101110110010101110001011100010100011101110111011100000111011101110111010001110110000101110111011101100001001000000010010001110111011100010110010001010111011101110111011101110111011100010111011101110011010001000111010101110111000001110001011101110101011100100111010101110110000000100111011101110100011101010111000100100111011001110111010101000011011100100111011101110010010001110100010101110111000000100111001101110111001000010111011101000000011101010111011101110011011101110111011101110111",
		"01110111011101110011011101110101010001000111011101100010000001110110011100110100011101110111011101110111011101110110011001110111011101110111000101110100000000100111000001100110011101110011011100110100011100010111001001110110011101110010010101110111000100010111010001110111011100100011011100100010011101110010011101000010000101000111001101110111011101100100011101110000011101110100011101110111011101110110001001100100011101110010010001110111001001110111000001110111011100010111011101110111011100010101011101010111",
		"01110011011101010111000001110111010101110111000001010100010001000111011100100010011101000100011100110111010001110001010101110111011101100111011100010010011101000111001101110000001101000111011101100111011101110111001101110101010001110010011100110111010001000110010101110101010001110111011101000111001101110111011101110111011101000111011100010110010001110001010101110111010100100111011101110111011100000001001101110000011100000111011101110100001001110111011101010111001001110111011101110001011101110111011101110111",
		"00110011011001110101011101110110011101110010011101110111010000000110010101100111000000010111011100000111000100110111001100010011011101110111000001110111000101110111010001110111000100110101011101110001011101110111000001110000000101110111011101110111011100100010011001100111010101100110011100100101011101110111011101110111011101110110011100110110011101000110000101110101011101110110010001110101000101010011011001110010011100000111011001110000010001110111011101000010000101110111011101110111011100100111001001000000",
		"01110100011101110111000001100111011101110111000001100111011101110111010001110011010001110111011101110111010001110111000101110010011101100111011101000111011101110010011101110111011101110011011101100111011101110011011100000110011101110001011101110110011101100111000101110111011101010111000100010010011101110111010001100111011101110111011101000111000001010111001000110111011100000010011101110111011100100010011100010111011101110110011100110111011100010111011101110111011100000111011101000010011100110111010001110110",
		"01110111011101110111011101100100011101100111011101110100011101110111011101100101011100010111011101000110011101110001000100000001011101110111011101110111001001100111001101110110001001110111000101000101011101110000000100100000000101000010011101110111010001110111011101110000001101000111011101110111011100100111011101000111011001110101011101110111010101110111011000010010011101110111011001000111011101110011011100000111011101110111011101110111000001110010011000010000000101110111011101110110011100110111011100100100",
		"01110111010000010111011000000000010001110111011001110111000001000111000100000001001001110111000100000111010101110111001100000111001101110111011101000111010001110101001000110010011101010111011101110010011101110101011100100111011101010011011101110001001001110111011101110111011101110101011100000011000100100101001101110111011100000111011101110110011101110100011101110111011100110001010001000011011101000110011101110111001101110010011101000111000101100110011101110111011101010110001101010111001101110001011101110111",
		"01110111000101000100011101110010011001000111011101110111010001110011011100010011001100100100000101100111000000110111000101110110010000000111010100100111000101000110011101110010010100100111011101110111010101110001001101110010001001000111001001110111011001110111001000010111011101110111000001110111011101110111011101110111010001110111011000010111011100000111010001110110011101010011010101110111011101110111011101110000011101100011011101110011011101110111011101110001011001010110011101010101011100000111000101110000",
		"00010010011101110001000001110111001100010111001000100001000001100111011101110001011101010011011101110111011100010111011101110000000001110111011100010001011101110111000101110010011101100100000000010101011001110111011101110111011101010101011101110111011101110101000001000011011101110001001001110111011101000111011101110111011101110010000000000111011101110110001101110110000001110111010101110111010001110111011101110111010001110000001100010111011101000101011100010011011100010111011100110100011101110111010001110111",
		"00100000011001000111010000110111011100100111011101110000001001010111011101110111010000100110000101000110011000010111011101010101011100010111010000010000001100000001011101110000011101100111011100000101011101110100011101110111011101110110011101000111000101110000010101110101011101110111011100110101010001000100010100100011011101000111000001110000010101110111011101010110011101110101001001110111011100000000011101110111011100100010011101010111011001110000011101110111001101110111011101110111010101000010011101110111",
		"01110110000001110001011100000111011100010101011101110010001001110011011101110000011101110001001000100111001000110100001101110111011101000111011101110111011101110111011101110100011101110110011101110100011101110111011100100010010101110111011101110111011101110111011101110001000101010001010001110011000101110011000100000111011101010111011101110100011101010010011101110111001001010111010001110111011101100010010100010111010000110110011101110000011100010110011101010111011101110101011100010111000001110111011101110100",
		"00110111000001110111011101010011000101110111001001110111001001110010011101110110010001110111011101110111000100100010011100100000010101010111011101110111011100000111001001110001011101110111010100010111001101000111011101110111011001110111011101110111011101000000011100100111011101100101011101110111011101110111001001110101011101110010000001110111000101110111011100110011011101110111011101000111011101110111011101010111011100110111011101110111011100110011001101010011011101110101011101110111000100110101011101110000",
		"00100111011101110111011101110111011101110111001100000111011101110010011100100111010100010100011100100111010101100000001000010000011100000111011001110010010000010111011101110111001001110111011000010111001100110111001100100111011000010111011100000111011001110101011101110100011101110110011101110010011101110111001100110100011101110111010000110111011101110110001101100110011101110111011100110111001100100110011101110001010101110001011101000111010000000111011101000111011100000111000101110111000101000111010101110000",
		"01110010011001110100000100010111011101110010011100000111011101110111011101010111011101100111010100000111001001110111011101110111011001110000011100110110011101110111010001110111000001110111000000010010000001000111011101110111011101110111010001110101000001110100011100010111011100010010011100110101011101110111011100110111011101110001011101110101011101110100011100100111011101110010000001110001010100000111011101110101011101100110011100100111011100110011011101000111011101110111011100000111011101110110011101110111",
		"01110010011101110111010001100111010101110001001101110111010100010111011101000111001101000000010001110000011100100111011100000111011100000111000001110111000001100111010101110110011101110101010101110010011101000110011101110111011100100010010000000011011101110111000100010111011101110111011101110111010001000111001101110111010000100111011101110111011100100010000000010111011101110000010001110111011101110110011101010111011100010010001001110111011101110111011101110111001001000000011101110001011101100010010101110100",
		"01110011011100010110001101000011011001110111011101000111011100000111011101010111011001000011011101110111011101110110011101110111001001100100001001110000010100110111000100010111010101110111001001110001011100110111011101110111000001110100011101110110011101110110010001110011011101000111011101110101001001000100010001110010010100000111000101110011011100110111011101000111010001110111011101110111000000110001011101110111011101110111011100010111011100010111011100010111011101110111011100000110010001110001000100100111",
		"00100100011101110111011101100111000000000000011101110111000001110010001100000010011100010000011001100111000101110111011101110111011101110111011101110010011101110010010101110111011101110111011100010111011101110111011101110111001100000111011101100111011100110111011101110111001000010111011100010000001001100001011100010111010001000001011101110111000001110111011101110001010100010111011101110111011101110111011101110111011101110111011101100111000000000111010001110111011100110111011101100010011001110111011100110011",
		"01110110011001110111011100110111011100010011011101010111001001110111011101110101011101110010011101110000011101110110000000000111001101010111011101100110000001110111011101110100011101100111011101110000011101100111001101110010011100010101001001110111011101110111011101110111001001110111011101110010011101110111011101110111011100000001011101110111001000010111001001110100001100100101010001110111011100100111011100110111011001110111011100110110011101100100011101110100011101000111011100100111011100110111000100000111",
		"01110111011001100100011101110101000100110111011101110101010101000001000001110000010001110111011101110111000001000011011101110111011101110111010001100111011101110000000100100111011101000000011100000011000000110011011101000111011101110111000001110111001001110100011100000111011101110111001001110111001001010010011101110011010101010001011101110111011100000101011101110111000000000111011101110111001000000101011101110111011001110111001001110111011100110111011101000111001100010111000001010100011101000010001001110101",
		"01110111011101110101011000110011001101110011011101100111010101100101011100000100011101110111011101110101000100010100011100010111001101110111011101110111011100100000011100000100001001100111001000110111011001000000010101010000011101010110000100100111011100110111011101110100001101110111011101110101011101110111011100110100001100100011011101110101011100000111011101110111011001100111011101010111010101110111010100010111011101110111000001110111011001110111000101110111011101010111010000100111011101010111011101000111",
		"00110111010000000111011101110111011101110111011101110111011101110111011100000011011001110110011101110001011100000111011001110101000101110110000100010111011101110000000101110000011101110110000001110110011101110100011101110010000101110111011101110011011001110111011101110010011101010000011101010000011101110101000101110000010001110111001001110111000101110011011101110110011101110000001001110111001101110111011101110100011101110111000001110111011101110001011101000000001000000011011100110111001001010111011101110001",
		"01000111010000010000011100100011010101110001010001110010010101000110011100100111011101110111011101110111000101110100011101110111011101010111011101110010011101110111011101100101000001110101001100010111011101010111000101110010001000010011011100010111000101110111011001000111011101110111011101110111000101110111011100010010001001110010000101110111001101110111011100110111010101110010011001110000011101110010011101110000011101110001011101010111010001110110001001100000000101110110011100110110000001110111010000010100",
		"01110111011101110111010000110111000101110010011100100111011101110000011001110111001100010111011100010111011101110111011100110111010101110111001001110110011101010101011100100011011101110111011100000101000101000111011101110011011001000101000001110111011101110111011100100111011100000100011101110100011101110111011101100111011101110111011101110001011101110111001001110111000101110111011100010111001001110001011101110111000000100001011101000011011101100111010001110001011001110111011100100111011101000111011101110110",
		"01110110011101110111011100100101001001110111010000100111011101110111011100100111011101110011011100010111011100100110001101110111001000110011011101110000011100000101001001110111011101110111011101110111010001110001011101110111010101100111011101110111011101110011011101010100001101110111011101110111011101110111010101010111011101100111011101000010011101110111010100100101000000000111000001110111000101110111011101110100011101110101011101110010011101110111011101110111000101000111011101110110001001110111011101100111",
		"01000000011101110011011101110001011100010111011101110000001001110001011101110111011101110111001001110111011000100011000101110000010101110010011100010111011100100111011101100111000001110000011000100111011101110011011101010111001001110111001000010111000101110010011101110111001100000111011101110110010101110001011101110001011101110111011101110111001001110001010100010111011101110111010001110111011101110010011101000111011101110001001101110111011101110110010001110110011101110111011101110111011100110111011101110111",
		"01110101011101000111001101110111011101110111011100100111011101110111011101110111011101110111000101110111011000010111011101110010011101110101001101110111001001110110000001110110010100000101011101110111010101110000011101110000000100000010011100100111000001110111010001110010011101110001000101110111011001010101000001110111001001010111011001110000011101110011000101110011001001000111011101110111000001110111011101000001010101110111010100100011011101110000011100110101011101110100011101110111011101110111011100000111",
		"00000111011000100001011101110111000100110010000000000111011001100000011101000111011001110111000101100111000001110000011101110111000000100111011101000100010001110111011100000100011001110100000101110101010101110111011101010111011101110111011101000000001101000100011100110000011101110111011100000010000001110011011101110111011101110110011101110001010001110111001101110011000101110111011100010111010001110111010000000011010100110111011101110111010101010011001101110111000101110100011101100111011101110111011101110000",
		"00000100011101110111011101010101011101100111001001110111011101110111011101110111011101100101011101110101011101110111011100010111011101110111011101110111001001110111011101110111011101110010000101110100011001000111000001100111011100110111011101100001000001110111011100100111000101110111011100100001011101110110011100100111001101000111011101110010000100010111001100010110011101110111011100110111011101110111011101110111000000110111011001110111011101100111011101010111000100110010011101110111011101010011011101010111",
		"01010011001000010100011101110100010000100111001001110111010001000111011101110111001000100111001001110110011101110111001001100010001101110111010001110111010101110111011101110010011101010000011101110101001101010101011100010001011101110010010001000101000001110111011101110110001101100111001100110111011101110000011101110111011100100111011101100111000001110100011101000111010001110111011101110011011101000001011101110111011100100111001001100111010001110111001101110111010001100111011101110111011101000111010101000111",
		"01110101011101110011000100110000000101110111011100010111010101110111011101010111011100010111011101000101001001110000011101110111011001110111000101110111011101110111011101110110010101110111011101110010011100110111011101110111011101000111011101110111000000110111001101110111001101110111011100000110011101010110010001110000011000100001000101110000011000100110011101110101000101110111001101100110001101110111000001010111011101110111011101110111000001110111010001010011011100110101000001110011011101110100000001000111",
		"01110111011101110111000001100111011101010110011001000111011101110111011101110111011101110111011101010111011101110111011101110111010101110111011101010111011101110111011101010100000101110011001101110000011100000001011101100111010101110111011100110011010101100110011101000111011101110111010001010111000001110111011101110110001001110111001001000111011101110111011101110111010000110111011101000111011100110111011101110010011101110111010001110000011001100001011000100111011101110100011101110111000101110110011101110010",
		"01110001011100110010011101110010011001110100001101110111011001010111011101110010011100100001010101000111011101110110011101100011011101110111011101110111011100100111000100000111010101110000000001110111011100000001011101110111000101110111011101110101011101110111001101110100011000010000010001100111000101110111011101110011011101110111011100010111000001110111001101110111010101110100011101110011011101110000011101110010011100110010000000110000001101100100011101110111000001110111001000000111011101110111011101110000",
		"01110001011100100010011100110111000100100011011101010111011001110111011100110011011000010111000001110111011101110111011101110111011101110011010000000111011101110111011101010111011001110111011100100001011101110110000001100111001001110011010001110111011101010111011100000111011100100011001101000111000101110111000101110010011101110111000000010111011100110111000100000111000001110111011101110011001101110111010100100111011101110110010001110111010001110011011100000111001101110111011101000000011100100111011101110011",
		"00110110011101110111011100010011000000010001011101110111000001110111011101010111011101000010010100000111011100110111011101110111011101110101011101110111011101010010011101000111011101000010011100010111011100000000000101110111001100110110011101110111000001110111001100010001011101010111001101110111001101110101011101110001001001110011011101110001001000010111011101010111011100100101000100010111011101000001011101110011001000100111011101010110011101110111011100010111000100100101010101110111011101110000011101110001",
		"00110111011100100001000001110111000001110111010101000111001101110111011100010111000100100111011101110000011100100001011101110101011101110011011101110111011100100111011101000111001001110111011101110111011001110001011101100011010101110111011101110011011100010111011101110111011101110110011101110110011001000111011101110000011001110001010100000111000101010111011101100111001101110111010101110111000001000111010001110111011101110111011101110011011101110111011101100111001101110101000101000111010001110110011101110111",
		"01110111011100010101010000000111000001110001001001110100011101110111011101110111011101100111001101000111000101110100011100000111011100010111011101110101011101110100011101110110011101000111011101110110011101110111011101110000011101110111011101110111001000110111011101110111011101110111011001110011011101110111011100000111011101110110011101000111011101110010010101110111000001110111011101010010001101110111011101110111001101110100011101110110011101110101011100000111011000010111010100100111001101110111011100110111",
		"00010111011101110111011101110010011100100111011101110111011100110111001101000111001101110111000101110100011101110101011100100111011101110111010101110111011100000111011101110111000001110010000001110100011001010111011101000111000101010110011101110110011101110111000001110111011001110111000101010111011101010111011101110111000100000101011101110101011101000111011101110111011101110111011101100111000001110101011101110100010001110100001001110101011101000011011101110111010001110111011101110111011101100111011101110100",
		"01110111011101010111011101000111000100010111010000000111011101000111000001110111011101110011011100000100011100100111011101110111001001000001011101110111011101110111000001110111011101110111011101010100000001110000011101110111000101000101010001110110011101110111011101110111010100110111010101000111011101110110011101110111011101000001011101100111011101100111000001110111010101000111010001110111011101110110011101110111011101110001011101110100000001110111010001110100001101110000011000010111010101110000011100110111",
		"01110111000100100010011101100111001101110111011101010111011100100111011101110011011101110111011101000111011101100110011100110011011101110000011001110111011101110010011101110110001101110100001101110100011101000100011100110001011101110111010000100011011101110111011001110111011101110100010001010111000001100111011101110000011101110111000101000111001000100111010100100111011101010111010001000111011100000000000101110111000000010111011100110010011101110111011101110111011001110001000000000111001101110111011101110111",
		"01110001011101110111001101110011011101110100000000010111011101110111011101110000011100000111011100110111010000100100011101110111011101100100011101110111011001010111010000000111011101110001011101110111011101110011011101110111011101100111010101110101011101110111010001110111011100100111011101110110011001110110011101110111011101110111011101110111011101110111011101110111001101100111011101100111010100110111011101110111011101110011011101110011011101110111010101110111011101110111000101000100011101110111010101110111",
		"01110111001001010011010101110111011101100111011101110111011101110111011101110101011101110111011101110111011101010011011101110111011101000011011101110100011101110001011001000111011101110111011100110111010001010100011001110011001101000001010101110100001001110111000001110010011100000001000100100111011101110111010101110111011100010111000001000111011101110111011101110111011101110011011101110111011100000110010001110111011001110111011100100010011101110000011001110111011100010111000001110000000001110000011101110000",
		"01110111011101110111011101100101010000000000010001100111010101100111001100110000011100010111011101110101011101110010011101100111000001110111001101110111011101110110010001000110011101110000011101110111011101110111010001110111000101110111011101110000011100010001011100010100011101110111011101110111011101110111000001110001011101010111011101110111011101010011001001110111011101110100011100100100011100000101011101000100011101110111000001110100011101110111010101110011011101110001011101110000011101110111011100100000",
		"01110111000101110011011101110011011001110010011101110111011101110110010001110111000001110111001100110000001001100011010000000111010101110010011100010010011001100111011100010000011101100011011101110110010100110111000000100010011101110111001001100110010000010111010001110111011100010111011101110111011100000111000101110111010001010010011100100011000001110001010101110111011100100000011101110111011101110010001001110111011101110111011101100111000001110111011101110101011101110111010101110111011101110111011101110111",
		"01010110011101110111011101110111011001110111011101110001000001110111000100010111000101010111001101110111011100010101011100100111011100000111001101100100011101110110010001010111010100010011011101110100001101110111011100010111011101100110011101100100011101110100000100110111011101100001001000110101011101110011011101110111011101110111011101110111011101110111011101110111011101110100011101110110011101000000011100100111011100110111011101110011001000110111011100000010011100000111011101010100011101010111011101110101",
		"01010111011100000101011101110001000100100111001101010111011101010010001100010111011101110111011100000111011101100111011101110101011001110001011101110000011101110111011101110100011101110111011100010001001001110011011101110110011100000111010100110111000000110111011101110111011001110100010100110111011101110111010101000111011101110111011100000111001000010011011101100101011100010111011101110001011100110111011100110100011101110111010001000111001101010101000101110001011001110111011001110111011100100110011101110111",
		"00010000000001110000011101100010001101110111011101110111010101110111001000010111010100000111011100100111011101100100001101010111011101110111011101010011010001110100000001110011011101110101011101110111011000110111000101110111011100010110011100010111011101110111011100110010011101110111011100000111011101110110010000010111011101110111011001110001011000110001000100000111011101010111011101110111011101110111001001110111000100000111010101100111011100010111011100110111011101110001011101110100010000100010010000010110",
		"01100000011101110111011101110111011101110111011101100111011101110101010101110001010001110111010000110111001001000111011101100101011100010001001100110111011001000111011101010000011000000101000100000011000101110101011101110111011100100010001101110110011100110111011101110111011101110110001001110101011101110111011101000111001001110111010101110100011101110100001100110000010101100011011101110111001101010111011101100111011101110001011101110001011100100000011100110111011101010110011101110011011101010110000101110111",
		"01110110001001110111010001010111011101110111011001100010011101110010011101110111010101110101001001110111011101110111000101110001011101110001011101110100001001110001001101110111001101110111011101000111001001010111011101110011010101110010000101110111011101110100011101110010001001100111011101110011011101110111011101110101011101000111000000010010011101110111000101110111011101110111001000110010011101110111011100110111001101110110011101110111001101110000011100010111001001000111000001100111001000010111011101110111",
		"01110111000001110110000101110101011101110110000001110111010101010111011101110000001001110011001000110111011101010111010101000101011101110111011100000001000101100111011101010111011101110111011100000000011101110001010101000111000001010111011101110010011000100110010000000011011100100111011100010111010101000111011101110111011101110001011100110101011101110111011101110101001001110111011101100111001001100001011100000001011101110111001000000110011101100011011101110001010000010111011101110011011101110111010001110100",
		"01110101011100010001011101110111010101110111011101110000000001110100010001110111011101000111001001110111011101110111000101110001011101110110011101110110011101010010000000100111011101110001011101100100011101110111011101110111011101100001000101010111001101110110000101100111001100000111011101110110010101110111011101110111011101110111011101110011011101110001011101100111000101110111011101110111011001010111000101100111011000110111011101110111010001110111010101110011000001000000001001010101010001110000011100010110",
		"00100111011101110011000101110111011001110111010101110111011101110110001001110111000000100111011101100110011101000111011101110111000001110100011100010111010001110110001000010001011100000110011100000101000001110111011101110101001001010111011100100011010101110011011101110111011001010101000000110011011101000101011101110111010001110111010000100000011101110111011101110111000100100000011100010101000000000111011101110111000000100111011100100001011101110010011101110111010001110001011101110111010000100111001001110111",
		"01110111011101110111011101110111011101110010000001110111011100010000011101110111000101000111011101110111011101110111011101110011011100100111011101110000011001010111011101110111000101110101011101110111011100010111010101110111011100110111011001100111010101110110011101110111010100000000011101110100011101110010010001100111000001110111011100100010011101110111001101110001011100000111011000000111011101110111010100100111000001110110011101110111010001110010010001110111011101110111000100100111011101110110011101110000",
		"00010111011101110111001101110111010001110011010100000011011100010010011101110111011101110111011101110111011000110010011101110111011101110111001101110001011101110111001000110111011100000111011100000000011101110111010101110000011101000011011101110111011100010101011101110101011101110000011101110011001101000111011101110111001001110010011101110111011101100111010001000010000101110100011101110000011101010110011101000111011000000010011101110011011100100010011101110100011100010111011100110110011101110010011101110000",
		"01000100010100100111001101110110011101110111011101000111001101110111010101110001010001110111011101110111011100100011011101000111000001110100011101110000011101110111001101110101001001110000011100110100011101110111011100100111000100010111000000110111011101110111011100010010011101000111011101110111011101100111011101110111011101110111011101110111011001010011011101100101011101110111011101110111011101110101000101110111000001110111011101100111010101110111001001010111010101110111011100010010011101110111011101110101",
		"01110100011100110111011001110111011101000111001101110111000101110101001000100110010001110111011101110111010101110111011101110111011100010010011100000001011101110001011101110111001001110111000001110110011101010100011101100111011101110101011101110111011101110000001001110000010101000111001000110111011001110111011101110111011101100101011100100001011001110111011101000111000101110111011100110111011101100111011101000100011100110111011100100110011101100101011100010110011001000000011101110111001101000111011101110111",
		"01110111011101110100011101110100011001110011011101000000011001110001010101000111011101110111011001110011011100010111011100100010011100100111001101110110011000100000000001110000000001110111010001110100011001110001000001000000000001100111000001110011001101110111011101110001011000000111011101110000001000010111000001100101011101110000001101110001011101110111011100000111010001010111001000100001000101110111010000000000010001100111011100100100011100010111011101110011011101110111011101110111011101110000011101110011",
		"01110111011101110111011101110111010100000111011101010111011101110111011100010100000100110000011101110111010001010011010001110001011101000001011101110001011100010111010101110111011101110111011101110011011100110101011100110101011101110111011100110111000001010111011101010101011101110111011101010001011100110111011001010110011101110111011101110010011101110101011101110111011101110111011101110111011101110001011101110010011001110111011101110111011101010111011101110110001101110111000101000011001001110111000001110100",
		"00110111000001110111011100110111011001110111001101110000011100100110011100010011011101110010011101110111011101000111011101010001011101110011011100010111011101100111001100010010011101110111001001010111011101110111011101110111001000010111011001110110011001110001001001110001000000010000011100000111001000010010011101010011010101110100011101110100011101110111010100010111000001010111011101110001011101010101001101110111000001100010011100100001011101110110011101110100011101110011011101110011010101110110011101010100",
		"01110111000101010110011100100111011101110010011101110000011101000111011001110101010101010111011101110000011101110111011100100111000101110001010001110111011101010111000101110110011100010010000001110111011101100000011001000100011101110111000001110001011101110111011101110111011101110111011101110001000001010100000001110111011101000001011101110000011101110101001101110111010001100000000101110111011101000100011100010011010101110111011101100111011100110001011100010111000000100001010001110010011000100010001101110111",
		"01110111011100110011011000000111011101110111010001110101011001010000011100000111000101110111011001110111011101110111011101110111010001110111010101000110011001010011011101110100001001110111011101110110011101110111011000110111011101010111011101110001000001110111011001100111011101000000011101110110001100100010001001110111011101110010011101110100011101110111011101110001011100100111000100000111011101100000011100010111011101110111011100000111010101110011010101100000010101110000001101100111010000010111011100100101",
		"01110111010001100111001000100010011101110111011100000110011101110111000101110111011101000111011100010111001101110100011100100111011100000111011101000100000101110110010101100010010101110111011101110111000101110100010000110010011101110111001100000111011101110111011101110100011101100111000001010001011000010111001101010100011101110111011100010111010101110111010000110011011101110110010101110110011101010111011101110000011100100111011101110101010001010001011100110100011101110001011101110111001000110100011101100111",
		"01110111011100110111011101000111011101110111010001100111000000010111011101110111011100100111010101110111000001110001010001110010010101010101011100000111011101110110010101010101011100010100010101000111011101010001011101110111011100100111011101110101011100100110001001110101011101000100010101010101011101110111001000000110011001000111010001000101011001110111011101110111011101000111011100010111000001110100011101010100011101110111011101110111011001110110011101110111011000010110011101110111000101110010011101100111",
		"01110111011101000111011101110111011100100000011100000001000101110001011101110000001100010111011101110111000101000111001000010111001101100111011101000111011000010111001001110111011101110010011101110111011101110111011101010110011101110111010001110111010101110111011101100010001101110111011101100111010101100000011101110111011101110011011100110111000000000111011101110111001001110110001101110111011100100111011101000011011101010000011101110110001101110111011101110111011101110111011101100100011101110010000101110100",
		"01110100011100000100010101110111011101110111001101110111011101110110011101110100011101110110001001110111010001110111011101110011011101000110011100010111000101110111011101110111010101000010000101110111000001110110011100000101001001000111011101110111010000010000000101110111010001000111000101100001011101110111011101110111011101110101011001110111011000110111001001110100011101110111011100110101000101110101010001110111011101110111011101110111011000010111011001110010011101110111011101110111000101110111011101110111",
		"01010111000101110111011101110111010001110111011101110111011100100011011101010000000101110001011101110111011101000000011101110011011100000111010000000111001001010111010001110111010000100100001101110111010001000100001000110010001101110001011101110110011101000111011101110001010101110111011100110110011101110010011101110100011001100111011100000111001000110111011101110111011101110110011101110011011101100111011101110111011101000111011101100000000101010111011000000111011001110111011101100010011101110111001001110111",
		"01110111011101110111011001100111011101010011011001100111001101000111011100000010001001110111011001010101011101110111011101110111011101010101011101110111011100000111011101110111000101110000011100100100011101110111011101110111000101010111011100010111011001110111011101110111011101110111011000010011000101110111011101110111001100010101010000000010011101000111011101110110010001110111011101000111011100100111011101100111011100000110011101110111011001110001011100010110001101110111011101100101011101100100011000000111",
		"01110010010101000111011101100010001101110001011100110101010101100111011101110110010001110111001101110111010000000111011101110011010001110100000101100111011101100111010101110111011000000011011101110111010101010000000101110111011100110111011101110111011101110011011101110111000101110111011101110101011101100111011001110000011100110111011001010111011101110010000101110000001101110000011101110101011101000010011101010111011100010111011101110011011101110111011100110111001001110111011101000010011100010110011101110111",
		"01110010001101110111010001110111011001110111001001010111011101110100000101110011011001110111011001110001000000100001011101000111011101110110011101100111011101010111000001110101000100000111010001110111011101010111011101110111001100110010000001110111011100100000011101110010011101110110011101110111011101110101011101100001011101110111011101110000011101110111001101110011000000110010011100110111011100010001011101110111000101110111001100010100011100010101000101110010011101000111000001110111011101100111011101110111",
		"01110111011101110111000101110100011100100111010100110111011100110111010101110100001101110111011101110111011100110111001001110111011100110111001001110001011001110111011101110111011101100111011101000100011100010111011101110111011101110110010101100111010101110111011101110111011101110111010001100110000001110111011101110000011101010000011000000111011001110001011101110111011100010111011101110111011100000101011100100111000001110111011101110010010001110111011101110111011101000111011101110111011101100100011101110111",
		"01000111011100100111011101000000011101000111011001110111000001110100011001110111001101110000011101110111011101110110000101110111011000010111010101000111011101110111010001110111011101000000011101110000011101110111011101110100011101110111010101110011010001000010010101000111001101110111011001000111010101110111011101000000011001000111011101110111011101010011011101110111011101110111001100010011010000100011011100110100011101110000011101110111011101110111011001010111011101110111011101110111011100110111010001110111",
		"01110111000100000111001001000011011101110011010000000111001101110111011101110111011100110111010101100111011101110111011100110110011101000111011100000111010001110111011101110111011101110111011101110111001000000111010000100111011101110111001101110111000100100111000001110110001100110000011101110110011101000101000001110111011101110111011101110011011101110111011101110100011100100000011101010111000101110111011101110010011101110111000101110101011101110111000101110111001101110000011100110111011100010001000000100111",
		"01110100011101110111000100000111001001110011001101100111000101110100011101110111011001110011001101110001010100010100011101000111010100110100001001110011011001110111000101100100011101110100010100110010011101010000000001110111001101110110000001000111011101110111011101100101000101110100011101110111011101110111011001110111011101100111011100110111001001110111010001110100011101110010010100000110011101110010011100100111011101110111011000100100011101110111011101110001011101110010011101110111011001110111011101110111",
		"01110111011101010011011100100011001101010010011101110011011101010000011101110111011101110101011101110111011101100111001001000111011101110010011101110001011101110111010101110000001100000111000001110111000001110111011100110110011100010100011101110010010001100001010000110111000101110111011101110111011101000000011101110100001000010110011100100110010101110111011100110111011101110101000001010001011100100111010101110111011100010111011100010011011101110000011100110111011001110111000100010111001000100100000101110111",
		"01110111010100010010011101110111010101110111001100100110010101110100011100010101010101110111011100010111010000110010011101110001011100100111010000010111011101110101011101110010001001110111000001110110010001100111011100110111011101010111010000000111010101110111010000010011010101110001011101010111011000100000011100010010011100110110011101110111001000000110010101010111010101110111011001010011000001110111011100000111000001100000011101110110000101110111011101110111011100110111010001110000010101000111011101110111",
		"01110111011101110111011100110001011101110111001000010001001001110111011101110101011101000111000101010100001001110111000101000111011101110111001001110111001101110111000001100010000001100110011101110111010101110111011101110101011100110110001101110111010101000111011101110111011100110101011100000110011101110101000001110100011101110111011101100111011101110110011101110111011101110111010000000010011100010111000101110111011100110111011101110111011101110111000001010101011101010111011000010101011100100111001001110010",
		"00000111011000010111011101010010011100010111001101010100011100110111011101110111011100100111011101110111010001110111011101100111011101110010011101110111000001110101001000110111001101110111011101110111010001110010001000000101011101110111011101110100011000110111011101110111011001000111011101110111011001010010001001110111011100110111010001010000011101110111010101110111011100010000001101110111011101110110011101110100011100110001000101110111011101110111010101110111011101000111011101100111000001110111011101110101",
		"01110111011101110101011101010011011101110111011100010000001001110110011001110101010001100111000101100111010000000100011001110111010101100011000100000111000101110111011101110110011101100001011100010111000000110001011100000011000000100111011101110111011101110111011101110010001000010111011101110100010100110010011101100111010101110111011101110111011101110111011101110111010101110110011101110100011100100111011101110101011101110111010001110000010101110111011100000111000101110111011101110000000101100111011100000000",
		"01110100011101010111011000010111000001000111011101110111011001110111000001110001011101110111011100110110011101110000011101110111010001110011001101100111011101110101010101110111011101010111000001110111011101110110011100010111011100010110011100110001011101110011000101110000001001110111011101110111001101110111001001010110011101110111011101110100000000000111011100110111000100010000011101110111011100000111011001110111001101110101011000010101011100110111011100100111011101110111011100110111001001100111011100010010",
		"01100111011100000111000101110000000001110111011101110100011001110101011101110010000101010111011101110010000101110000010101010110001000110000000101110101010000100011000001110111011101100111001001110010001100110101011101110010011101100111001001110100010001110111001101110111011101110110011000000111011001110010011101110110001000000110010001100111011101100110011000100111011101110111011100010101001001110111011101010100000100000111011001000111011101110011001001110111010100010110011101110101011100010011011101110111",
		"01100111011101110101001001010111000001100111011101110111011101110010011101100111011101110110011101110111011100100111010101110010010001000101000000010110011101110111011101010010011100010010011101000110001101000000001101010111000101100100011101110101001101110111011100010111010101110100011001000001000101000111011101110011011101100011011101110010011101000011000101010000011100000111010100000010011101110111011100000111001000010111011101110111011101110110011101110111011001110100000101110111011101100111011100000000",
		"01110111011100000111011101110010011101000111010001110111011101110111011101100111010101110111011100010111011101000111011101110111011101110000011101110111011100000111010001110111000101110110011101110011011101110100010001110111010101110111010100000100011101110110011001000111011100110101011101110101011101100101011101110001011100110001011100000111001001110111010001100010011100100111001101110111011100000010011101110111011101110111011001110111011101110111011101100111011101110111011101110000001001110010000101110111",
		"01110111011101110111010101110101011100110111011101110100000001110001010001000111010101110101011101100111011101110000010001100111000101110110001001110010011101110111010001110010011101110101011100000010011101110111000001100111011101110111011100000001011101110111011101110111011100010011011101110001011101000111011001110111011100010111011101110111011101010000011001110101011101100111011100000101011101110111010100000111011101110101011001110111011101110010011001100111011101110111011100110100001001110011011101110010",
		"01110111011101110111010000000111011101110111000100000111011100000010011101110111001100000111001101100101011101010111011101110111000001110001011100100100011101110011000001110100011101100111011101110111010100010100000101110001011101110011000000110111010101110111010000000111011101110111011101010111010101110111011001110111001101010111011101010111011101110110011101000111011101110101001000010111011101110101001001110011011101110001011001110111000001110111011100000111011100010111010001110011001001010001011101010111",
		"01110001000001110111011101110110011101110001011001110010011101110000010001110001011101000111000001110001011001100111010101110111010101110111001101100111011101110001011101110111011101010111010101000111011000100111011101110111011100100000000001110000001101110111011100100111011101110111010000110111011000000111011100110111011001000001001000010111011101110111001000010111011101010111001001110111010101110011011101110110011101010010011101010101011101110001011101110111011101110101011001110111010001000111001101000111",
		"01110000000001110001011101100111011101110111011001110111011101110111011101110010011101110111011101110111011101110101011001110110010101110101011100100111000000100001010101110111001001110111000101110100011101010011011001110111011101110101011101110100011101100001011101110111011101110011011101110011011101110111001101110111011101110111011101110001011100100111000100100111011101110111010000100011000101110111000001110111011101110111011101110010010000110111011101110111000001110111000101110111011101110111011101110111",
		"01110111011100110101010101110111000101000111001001010111000001100001010000100111011101110111001001110111000101100111000101110010011101110110001001110100011101110011011000000111011100010111000101000101011101110111011101110111001101110101001101110111011101110111010100100111001001110111011101100111000101110100010001110001011101110111011101110111011101110111010100110100011101110010011001100111010001000111011101100111001001110111011101110111001100100111011101110000010001110010011101110111011101110010011101100111",
		"01110111011101110111011000010111001100100111010101110000001001110101001001100111010001110111011100110011011101110111001001110010000000000000011101010010011100110111011001110100001001110110010001110111001001100111001001110111001100110111010000100111001101110111001000010111011101010111011101000111011101110111011101110101011101110101001101100111000101000101011101110111011100100100000100000111011101110110011101110101011101110111011001110111011100100111011101110111010100000111001000000111010101110111000101110111",
		"01110100001001110100011100000111011101110111011101110001011101110111011101110001010000110111001000100111001000110101001101110010011100110111011101010101001101110110011100110000011101110111011100100111001101110111010001110111010101110111001000110111011101110101011101110111011100100000011001110100011101110110001101110001011100010011011101000111000101110010000101110111011101000111011101100101001101110111000001000001001000100111011101010010011001110100000001110010011100100101011101000111010101100101011101010111",
		"00000111011101100111011101110001011101110000001001110111011101110111011100000010011101100001011100110111011101100111011101110111010001110111001101100110011100000111011101110001011101110111011100010111011001100111000100010111011001110111011101110010011101110111011101110111011101110111000101110110011101110101001000010111011101010111011101110110011101110111001100100011011101000111001000110111011101110100011100000111011101110111011101000111011101110111001100100110011101110111011101010000011101110100011100010000",
		"01110111011100110111010000110111010101110111001000110111001001110111010001100111011000100111011101110111011101110110011001110100011001110001011100100111011101110101010100100111011101110111011100010111000000110110011101110111011101110101011100100010011101110111011101110111010001110110001101010111011101110111011101100111010100110011011101000101000000000110011101100011000001100101000100010111011101110111011101110010001001110101011100010011011101110000011101110111011101110001000001110111000101110111000101110111",
		"00100010011101100111011101110111011101110111000101110111011100100000011101110100011101110111011101100111000101110000010101110000000101110111011100100100000001110101011101110101011101010000011101110111011101110111011101110010011100110100001001110000011101110010011101110111001000010111011101110111011100110100011000110111011101110110001001110000011101110101011100000101011101110000001101000111011101110111011101000111011101110111001001000101011001110111000000000011000101100111011101110101001101100000000101110111",
		"01100110010001010110011101110001011100110011011000000110000101110000011101110111000101110111000100100011010101100111011100000111010000000010011101110111011101110001011101110111011101110100011100000111011101110000011101110111011101110001011001100111010100100000000001110100011101110111010100010111010101110010011101110100011101000001011100010001011100100110011101110101010101110111011101110000001000110111011100100111010000010111010001000111000000110111011101000101011101110111011101110111011100100010011101110001",
		"01110110010001010100011001110011011101110001011101110001011101010110011101110000011001110101011101000111011101110010011101110100010000100101001000100100011101110100001000100000000001110111011100010111011100000001011100110111011101110010011101110111000000100101000001100111011001010111011101110111000001000001011100010111000001000111011101110000011100000001011101100011010101110111000001000111010101110111011100000111011101110111011101110010011100100000011100010111011101110111011101110111010001000111011001110111",
		"00000000011001110101011101110111011101010100011001100100011101000111011101110101010001110111011101110101011101110111010101110111011101100111000100100111000101110011011000000100010101110111000101110111011101110111010001110111011101110111011101110111011100110010011001000111011101110101011101110111011100000111011101110111011101110100011101110111010101100011011101110111011101010111011100110111011101110000010101010110011101110000011101000111010101110111011101110111010001100011011101110111011100100111011101100000",
		"01110000011101110111011101110111001101110111011101110000011100010111011100000111011101000100011001110111011101010100011101000111001101110111011101010100011101110111001101110111010001110111000101110110010101010111010000000111011101110111011100100111011100010111010001010111011100100111000101110111011101110111010100100111010000110101011101110111010101010111010000010111010101100111011100110111011101110001000101110111010100100111010100100010011101110111010101110001011101110111000101110000000100000111001001110111",
		"00100111011101100111011101100011000001110111000100100111011101110111011101110100011100000111000100010000001001110101011101010111011101110111010000110110000101010111011101110111010001010101011100100111001101000010011101110111011101110001010101010111010101110101011101110111011100110000001101110111011101010111011001110111001000000111000000100111001101110111011000010000011101110011011001110101011100110000011101110111001001110001011100110111011101100111010000010010001001110111010101110111011101110111010001110111",
		"00000111011101110111011101110111001000000111011100110111000001110111010001110111011100010010011101110111001000100111011100110110010001110111011100110111011101010110011001000111011101110000011100110111011101110111011101100110011101110111011101110110011101110111010101110111001001110111001001010000001100110111011101110011001001110111011101100011011101000100011101110111011101110111011101000101011001110001010001110001001101000100011100000001011101110111011101110111011101110111011101110100011101110011001101100011",
		"01110101010101110111010001110111001001110111010101110111010001100111000001110111011101110111011100100011000000000111011001010100011101110011011101110100010001110111011101110001000101110100011100000111000000100111011100010111000000110101011100100111011101000111011100000111011101110111011101000111000001010011000101110110000000000000011001110111000001110111011101110111011101110000011100010111011100010100011101110111011101110111011101110110011001110001011101000111011101110111011101110111011101000101011101110000",
		"01110001011101110111001100010101011100000100011101110111001100010111010001110111011100000011011101100010011101110110000000000111001000000000001101110111011100000111011001110000000100100111011100000111011100000110010000010111011101000001011101110111011101110111011101110000011100110111011100000111001100010010010101100111010000100101011100010111011101110000000101000110011101100111001100000111011101000001000001110111001000100001000001110010001101010110000100000001011101110101011101110111011001110000000101110111",
		"01110111000101100111011101000111001001110100011101110000000100000100011101110001000001110100001101110111000001110111011101110100011101110111000000100010011101010110011101010111011001110111000001110111001101110011010001110110000101110001011001110110011001110110011001110111011101110000011101100001011101010111011101010111011100000111011101110001011100000111000101000110010101110111000001110001010101110111011101110101011101110001011101110111011101100111011100010110001000100111000101110111011101110111011100010111",
		"01110111010101110010011100110111000101110111011101000111011101110111010000010011011100110111001001110111000101110111011101000001011100100010001100000110001100010111000000100111010000100111011101110111011101100111010101110000000101010010011101110111011101000111001101110111011101000011011101110011011001100110000101110010001001110111011101110101011101110001011101000101001101110011011101110101000001000111011101110111001101110010000001110111011101110010011101110011011101100111001100010111011101100101011100010001",
		"01110111011101000110001000100010001101110101011101110111011101100111011101110111011101110111000101110000000101110010011101000100011000000111001000100111011100110000011101100101011101110111011101000111011101110111001101110001010000110111000001110111011101110110011101110101011101110100010101110111010100000111011001000111000001110010001101110111011100110011011101000000011101110111010101100111010000000001011101100111011001110110011101110001010001010111011101110111010100100111011001110010011100000111011101110111",
		"01000111011100100111011101110100011101110010011101110001011101100111011100110110000001110010011100110111011101110111010001110111011101110000011101110111010101110001011101110010011101110111011101110111001001110111011101110111011100010010001001110110011001110110011101110001000101110111011001110110010001110111000101110011011101110000011101110111011100100111010101110111011101110111000001000111001101110011011101110110011101110111011101010111001101110100001100010101001001110110001000110111010101110111011100000010",
		"00010111011100000111010100000111011001110111011100100110011100110111010100100010011100110111010100110011001101110000001001100110011100010111000001110111000100100101011101110000001001010111011100000000010001110011011100110010011001110111011100110000011100100111000000110011011101110111011101110111011101110111011100010001011101110101000101110111011101110001001101110001011101000111000101110111010001110111000001110111010101110111000100110111011101110111010101000110001001010000010000100101011101110111011101110111",
		"01110011001101000110001101110101010001110111011101110111011001110111011101110111000101110001001000110111011101110000000100100111011101110111011101110111011101110001011101110111000001110100001001000111001001110000000001110111011001110010001001110111010000110111011001110101011101100111010101110111011100100111011101000100010000010111011101110111011000010010010100100011011101110111001000100111011001110111010001110000011101110111010101010110000001100010011101110110010101110010011100000110011101000000000101110111",
		"01110111011100010111011100100111011000110110011101110111011100100111010101110110000101010010000101110001010001110111001000010010001001110001011001110111011101110111011100010111011101100111010001110001011100110111011101110111011100000111011100100000011101110000011101110111011101110111011101100111010001110111011101100111011100010100011101110000011101110111000001100011011101110110010001110001011101110111000001100111011101100111000101110111011101110110011101110100001101110111001101110111001101110111011101100111",
		"01110111011101110100011100110111001001110011010001110011011101110101010001010111011101110111011101110111011101110011011101110001011101110001010001110111011000010001011101110111000000100111011101110111010100100111011100110111011001110111011101100111010001000001011101110011010101110111011101110111011100100111011001110111011101110111000101110111010101110111011101110111010101000000011101110111011100110001001001110111001001110010001101110010011101110111000001110110001101110100000000010110010101110111001101110111",
		"00000110000100010001011001110111000000110111011101110000001000000011011001100111010001110000011101110001001101110111000001110011000001110010011101110111010100000111011101110101000101110111011101110110011101110110011100000001011101010000000001110111011101110101011101100111011101110001011101110111001101110101011101000111010001110111011101110010011101000111010101110000011101110111011101110111011101110111001101110011000000000111011101110000001101110100011101110111010100100110011101110111011001100111011100100111",
		"01000111011101110111001001110111010001110110011101100111011101110111011100110001011101100100000001110111011100000101011100110111011101100010011101110111001000000111011100110100001100110111001101100001011101110100011001110111011101110111011100100110001001110111011101110011010101100111011101110101011101110010011101000110001101110111010001000111000001110111010101110111011101110111011101110101000001110111001101000110011101110011011101010101010001110111001100100111011100100111011100110010011100110001000001110111",
		"01110111001000010011000001110101011101110111011001110111011101110111011101100111000001110111011100000111000001110111010000010111011101000001011101000111011101100111000001110111011101100111011101110100011000110111011100010111011101000100000101110100011101110111011101110101010101010111011101110111001000100111010101110010011101110111001000000111011101110111011000000111011101110101011100110111010101110111011101010111011101110101011101110000000001110110011100000010000100100111010101110111010101000111011101010011",
		"01110010011101000111011100100111011101110111001001000100011101110111001101110110011101110111011100010111010001110111010101000001000001110000011100100000011101100011000000010111011100100111011100110110001101110111011101110111011100010111011101110000011100100111011101110111011100000111011001000111011100110011011100000111011101100100001001110011011101110011011100110100000000110100010101110111011101010010000101110111000101110111011101010111011101110111011101110111000000100110000100100111011100010011011100010010",
		"01000100011101110000011001110111011101110101011100100111011101110111011101000111011101110111010001110010011100010111001101110101011001110111011101110111011000010111011101110111010001110111001101110111011101110111000100100010001100110101000001110100011001110110011001110111011101110000011101010000011101110111001001110000011100100111011101110111001001110001011101100111011101110111010001110111011100100001011101110111000001110110011100010001011101100100011101110111011101110111011101110111010101110111011101110101",
		"01000111011001010100011101110101011000100011011101110111011100000111010001110110011101000111011100010111010001110111011100000111011101110110001001110111011001110111011001010111011100000111010101110101011101000111000001110101011000110110001101000111011101110111011101110111000000110101011101110111011101010011011101110111011100010111011101110010011101010011011101110011010001110111000101000001011101110011011101110100011101110111000001100001010101110001011101110000011101110111011101010011010001110000011101000111",
		"00100111011101110111011100000111011101110111011100100011000100000111001001110111011101110111011101010111001101110000011101110111000001110111010101110111001101110010011101000001011101110111011101110111011100100111011001110111010101110111010001110111011101110111011100100111010001110000000001110011011101110111011101110100011101110110000001110011011101110110011101110010011001100101011101110101011101110000000001000111011001110111001001010111011101110011011100010100001001010000011101010111011101000111010101110111",
		"00000111010101110111011001110111011001110111011101110111010001110111011100110110011100110111010001000111011100010010000001010111001101100111000001110000011101110111000101110111011101010111011100110101000101110111010000110111011100000111011101110111011100000111010100110110011001110111011001000101011101110110011101110101011001110111001001000010011100000111011101110111011101110111010000110111001101010111011100110111001000000100011101110111011100100111011101110010011101100111011001110111011101110111011101000000",
		"01010111001001110111011101110111011101110111011101110111000101000111011101110111000101110000000101110010011101010111011101110011010101000111011101110111011100100101001001110111000001000111011101100111011101110111011101110101000101110111011100110111000001000010011101110111011101100111010101010010011101110111010001110001010101110111011101110111000001110111011101110111011001010001011100100111011101110111011101010010010000110111011101110010010101110011001001010011011101010111011101110101011100110110011101110111",
		"01110111011101110111011101110110011101110001000001000011011101110100010101000110001101110111011100010110011101110100000001100101001101010110011100110111011101110100001101110010011101110111010101110101000101110110011101110011011101110111011101110100000101010111010000010000001000100111011101110111011101110111001001110000011101110111000101110111000001110111011101100100000100110101011101110111010001110111011101110011000001010101011101110000011101110101011100100111010100100111011101110111001101110111011101110111",
		"01010100011101110110011101110000000101010011000101110101011101110001011001110011011101110110011101110111000101100110011001110111010001110001010000100111011101110111011101110010010001110111000100100111011101010010000101110011010000110111011101110000011001110001011101110010001000110111001001010100011101110010011101110101011101110111001001110111011001010000011100010000011101110000010101110111010100000011011101000111010101110111011101100011011101110111011101010111011101110110011100000111011101010011011101100010",
		"01110111011101110101010101010111011101100010011101110101001100100000011101110101010101110011011000010111011100010101011101110111011101110111011100000111011101110111011101110111011001100101011101110111011101110111011100100111000001110000011101110000011101110111011100000111011101000111000101110001011101000111011101110111011101000110011101110000010001110110011101110111011100010000011101110111000101110111011101110101011101110111011101110111011000100111011101100000001000010111000101110111011100100000011101110110",
		"01010111011101110101011101000111011101010111011101110111011100010111001001010101011101010111011101110011001001110100001001110001011101110001011100000101011001000111001101110111010001000111011101110111000101100001001101110111011101110111001001110111011101110100011101110111011100010110011101000111011100110111011101000001000101110011011101110001011101110111011100000100011101110111011100100000011101010111011101110111010001100110000000110110001101110111011101100111011101110111011101110111011101110111011100000011",
		"01110100001001000010011101110000011101110111011100000111001101110101011101110101011101110111001001110000011101010111011101110111011101000111011100000111011000010111001001100010011101110001011101110111011100000111011101110111000000100100011101110111011101110101000000110111010101110111011101110101011100110111011101110011010101110111010101110111011101110110011001110111011100110110010001110111010101110110011101110111010101110111001000110111000001110111011000100110011101110011010001110111011101110111010101110111",
		"01110010000101110111011101110010011101110111011101110111011101110011010000100111011101000111011101110111011101110011000001110010000100010111011101000010011101110111001001110000000100000111011100100111011101110101011101110111011101110110011101110111001001110001000101110111011101110000000001110100011101110111000001110111001001110111011101110110011101110111011100000110011101110111011100010111010001110111000001110111011101110110000100110100011100100010011101110111011101100001000001010111011101010010011101110111",
		"00010111011001110111011101110111011101000010001001110111011100110101001001000111011101110011011101100111001101110111011101110100001000110111010001110110011101110111001101100100000101010001000000000001001001110101011101110111011101110000011100110111000101110111010001110000011101010111010101110001011101110010000101110110010101010111010000000111011001010111000100010100001101110010011101110111011001110100011101110101011101110111001100010001011101110111011100100111001101110110011101110100011101110001011001110011",
		"01000111000100100111011100000111011001110111010101010111011001010100011101110111010001110010011100100111011101110010011000000010000101110111011101110110011101110111011101110111011101000111001101110100011101110111011101110000011101110010001000010000010101110100000000110001010000010100011001110111011101110110011100010110000100000111011100000101011101100111011101100111011100010111010100000111011101110110011100110111010001010001000000000111011100010111011101100111000001000111001100110111011101110111001101110000",
		"00100010010001110100010001110111011100000111001001100111011001100111011101110111011101110111001101110111011101100111010101000111001101110111010101110010011101110111000101110111000101110111001101110101001101110111000101110011011101110010011100010001011101110111011100010111011101110100011100000001010101110010011001110101011101100111011101110001010001110100010001110111011100110000001001010111000100010110011101110010011101110111011101110111011101110101011101110111011101110111011101110011010100010111001001110100",
		"01110101001101110100011100010111011100110100010101110111011101110100011001110101011101110100011100100111011101110011011101110101011101110111011100000111011100010101001101110100001101110111010001110111011101110111011101110111000101110111010001110111011101000111011100000010010001110101011101010111011101110010000101110010011100010111010101110111010101110111011101110111011101110010011101000111011000000101011100010111011101000111001000010111010001110111011101110111011101110111011101110111011101110111000101000111",
		"01110111011101110110001000100110011101110111011101110011000101110100011101110111011101110111010001110101011101110111011100010111001001010111001000000111011101110111011101110010011101010010000000010111000001110101011101100000011101110111010001110111011101110001011101110010011101110011010001110001011101110111011101110110000000100111011101110111011100100010011101110111011101110111011101110111011001110011010001110111011101110011011101110101001100110111010001110111011100000111011101110111000101110011011101110111",
		"01110001010101010010011101110100011100000111001001000100011100010011011101010011011101110111011101110110011100000010011000110111011101110011011101110111001101110111011101110101011100100001010000100110011101110001011101000011011101110111011101110000001100100010011101000010010101110100011001010001011101010000010001110011001001010010010100000111011101110100011100010111011101110101011101110011011001110111010101110101001001110101010100000000011101010111011001110100011100000010001101110101011100100011011101110111",
		"01010111010001110111000001110111000100010110001101110111001101110111011101110111011100000101011101110010001101110111001101110110010001110111011101110111011101110111011101010010001101110100000101110111011100000111011101110011011101010001010100000111011101110100001001110110011001110111000101100111011101110000011101010110011101110111010001110111010001110011001001110111010001000111010001110111011101110110011101100111011101110111011101110111011101110111011101110111011101110111001001010101011101110111011100010111",
		"00100111011100010111011101110111011101110111010000000111011100110010011101110011001001110111011101110100001000010001011100100101010000000011011001110111011000000111011101110001010001110111000101010100011101110000011101110111001101100111011101110101011101110111010001110101000101110111010001110111000001100111011100110111011101110111011101110111011001110100000101100100011101000111000101110100001001110111011001110100011101000111010100010110010001110111001001110111011101110111010101110111011001110111011101110011",
		"01110111011100110111010000110011011000010111011101110111011101010111011101100000011101110111011100110111011101000111001000110001001101110111000001000111000001100010011101110110011101110011011001100101000101100111001101110111001101110000000101110110010101110111011101010001000101110101011101110101011101110111011101110111011100110001001101110111010100010111011100100011011001000101011101010111011101110001001001110101010001110001001000010100011101110100011101010111011101110111001100000111001100110111001101110111",
		"01110010011101110101011100010000000000110111011101100110011101110000001101110111011100100100011001110010011101110100000100000111010101010111011101110101011101110111011101110111010101110111011101110000010001100111010101110111011101010101011101110111001101110100011101110111000001000111000101110111011101110110010101110010011101110100011101110111000100000010001101000111000001110011011101110111011101100111011100100111011000010011000001110111001001110111011101110000011101010111000000010111011101110111011101110011",
		"00010110011101010111010101110111001100100111010001110111010001110110000000000011011101010111000101110111000001110111011101110111000101110100011101100111001000110111000001110111011101110111001000110111011100000111011100100011010101110000011101000000011101110111011101000000011101110010011101110111011101110111000100100111011101110101011100110111011101110000000001110010011101110111011101000111011101110111011101010111011101110111011101010100011101110000011101110111011101010010011101110111011100100110001001110111",
		"01110000011101000010011100010111010001110111011100100111000101110111010001110111011100010111000100000100011101110100011101110001011101110111011101110111000101100111011101110111010101110111011101010111000101110110011100100001011101110101000000000111010000010111011101110100010001000110011101110000011101110111011101110111001101110111011101110111011101110111000101110111011001110111011100100111000001110110000101100111011101110111011101110101001101110111001000000111011101000001011100000111011101110111000001110001",
		"00000110011101110111011101110010011101110111011100110111011101110110001001110111001100100111011100110111010001110111011101110000000100100011011001000111011101110111011101110111011101110000011100000111011101110111011101000011011101110011011100110111011101110111001001010111011101110111011100010111011101110111011101000111011100010110001000010000011101000111011101110010011101100111001101110011011101110110011101110010011100000111011101110111011101010111011101110011010101110111011101010111011100110100011101110111",
		"00100010011101110111011101110111001001110111011100010111011101000101010000110101001100000011001100110000011101110100010001100001011101110111011001110110011100110001010001110110011101110101010001110111000101110111001101110111011101110111011101110110011101110111000101110101011100010100011100000111010101110111011000010101011100100100011101110111010101110011011100110001010000000111010001110100001101110100011101110111010101100111011101000011011101110010011100110111011100000111010101110111011101110111000001110111",
		"01010111011101100001011101110111000001110111011101100111001000100111000101110111011101110001011001110111011101110111011101110111011101110111001101110111011101110111011101100111011100000001011101110111000001110111010000000001011101110001010001110011011100010111001101110000011100010011011101110010011100000111011101000001011101110111011101110111011101110000001101110000000101110010011101000001011101110111011101100111011101110111000101110010011101110010001000100100000101000111011101110111011101100101011101110111",
		"01110101000101110010000101100111011101010100011101010111011001110111011101110110010001110111010000110101011101110111001001100011010001100110001001010111011001110111011101110111011001010100011101110111011101110001010101110100011001110001010101110100001101100111011100000001011101110111011100110100011101110111011101110111000101110111011100110010011001010111011100100101010001010101011101110111011101110111011101110110011101100111000101110111001101100111000101000111001101110111011101110001011101110111011101110000",
		"01110010001000110111000101110100000001100110010101110011011100010111010100000111001001010011000101110010011101110100010101110111010101110111001000110110011100100111011101110110011001110011010001110100011101110111011001000000010000000100001100100010011101110111000101100111000001010111011100110110011101110111001001000110000101010011001101110100011001110110010101000111001001110111010101110111010001000101011101000111011100000010011101110111011100010111011100110001011001110111011101100111011100100010011101110111",
		"00000111011101110111001101100111011100010111011101110111011101110111011100000011011101000010000101110011011101110111010000100110011101110111011101110011011100100011010101010100011001110111000101110111011101110001011101110111001101110010011101110011011100010111011101110001001001110111011101110111011101110100011100010111001001110111011101110000011101110011011101110111011100010010010101110100011101000111011100110111011100000110011100010111011001100010011101110111001101110111000101110111011100110011000101110111",
		"01110101011101010100011000110111000001110111011101100110011101110111011100110111011101110010011101110111011101010111011100100111011101110110011100110111011101100010011101110110011101110111011101110001000001110111011101110011011101100111011101110111010001000111011101000111011101100111000000000010001000100111011101100110011100100011010101110110000001100111011101000110011101110100011101110011011101110111011100100110011101110001011101110111011100110011000100000111011101110111011000100111010101110001010101110111",
		"00110110011101110010001100010000000000110101010101110111011101100100010100000111011101110111011101110111010001110111011100000111011101110111010001110100010001000111000100110111000001110010000000100111011101110111011101110100011101110011011000010010010101110111011100110111011001100100001101010111001001110111000001110100011101110111001001110001011100100010011101110101011000010001011100010111011101100111011101110111011100100111001001110111011101110111011001110110011101100111011101110111011100010111001000100001",
		"01000011011000000111001001110011011001110000011100000100000101010111000001110010011100110111011101110001011101110111011100000101011101110011011100100011011101110111011101000000011101010101000101010111011100110111011101110111011101110111011101010100010100100110011101110111011101110111011101010000001001010111011001110111011101110101001001110001011100000011011101000100010101000101011100100111000001110111000100010001011101110111011101100100011101010111011100100101011101110000010001000111011101110101011101110110",
		"01110111011101110111011101110010011101110111010001110111010000000101001100000111011100000010011101000110011101110111011101100101011101110111011101110111001101110111000100000001011101110111000001100111011101110110011101100111001101110111000001110010011101000111000001110001011100110000011101110111010001110111001100010011011001010001011100110000011101110000010000000111011100000001001101110111000101110110001001110010011101110111011101110100011100000111011100110000011101000110011100110111011101110111011101110111",
		"01000111001100000111011101110110011100110100011001110001011100010111001101110101011101110111000001010000000000010111011101110110011101110010010101110111000101110001010001110100010101110111011101110111011101110100011001110110001101110111000101010111011101100111011101110011011100110101000101110111001000000111010001110111010101110111010101110111011001110111001001110011011101110111011101110110011100110101000101110111011101110100011101110111011001110111000101110000011101110111011101110111010000010100011100010111",
		"01110000000001100111011101110110011101000100011001110110011101110111000001110100011001110111001001000110011101110111011101110111011001110111010101110111011101110000010001110111010101110111011101110011011100110101000001110111000000000110011101110101001001110010011101000111000101110111010101000111011101110111001100010011011101110111010101110111000001110100000101000111011100100111011101110111010101110111011101110111000001110110011101110111011100100100011100010111011101010111000000100111011100010111011101110100",
		"01110111011100110111011101000111001101110111010100110111011100000111011101110110001101010111011101110111011101110111000001110111010101110110011101000110010100110001011100000110011001110000011101010111010100000010001001010111011101110111001001110111011001000111011101110110011000100111011101010111011101110111000001110111010001010001011000100111011101110011011101100000011101110111010001110111010000010111011101110111010100000000000001110001011101110111011101110111000001110111011101110010011101110111001101110101",
		"01000111011101110100011101110000001101110111001000100010011001110100011100010111001001110111000101110110010001110001011101110111010001110100011101110111011100110111001000100101010001110111011001110111011101110101000101110111000101110001011100010101011101110000011101110001010001110101000101110000011100110111011101100011011101110111011101110110011101110110011100110001010101110111011101110011010001110111011101110011011001110111011101110110011101110111010101110111011101110001011101110111011101110110011001110110",
		"01110111011100000010000101110011011101110111001001110101011100000111010100100111001001110100011101110111011101000011000001110000000001000001000101110100011101110101001100110111011100000111011101110111011101110111011101100111001100110111000101110111011101110110000100100011011101110100011100000101011101110111010101110101011101010011011101110111011101110100011100100011001100110100000100010111001001100011011101110111011101010111011101000111000000000011011100110111011101110010001001110101000001110011011101110110",
		"01110111011100110010011101110111011100000111001100100010000101010111001001110010010101110110011101110110011101110010011101110111001101110111011101110011011101110110011101010011011101110000011101110011011101100101001001000111011101110111011100010111001101110111011101000000011101100010000101110101011100110010011100010011011101110100001100110011011101000111010101110110011101110111010001110111011101110000010001110001000001110111011101110111011101110111000101000111010001110111011101110101000001000110000001110111",
		"00100111011101110111011101110001010100010111010101110111011101110111011101110111000001110101011100010011000101110101011100110100011101110111011101110001011101000000010101100111011101110111001001110011011101110111011100100010011101110001011100110101001101110111001001110001011101100100011101100011001101110111010100100011011101110010011101110111001101110111000101000001011001110111000101110111011100100111011100110111011100010110011100100111011101110111011101110111001100110111011101000111011100010111011101110000",
		"01110111011101110111011101110111000101100110011101110111011100000111011101000111001101110111001101000111011100010111011100010111010101110100011101110000001101110011011101010111011101100111011100000111011101110111011101110111010001000111011101110111010001110101010101110111011101110111011100100010011101100101011001110100001001110111011100100000011101000111011001110000011100000011011101110111001100000001000001110111011101110000010101000110011100100000001101000101000000000111011100100111011101110010011101110111",
		"01110111000001110111001000110001011101110111010001110000000101000111011101110101011001110111001100000111001001110111011100100000010101110111011101000110011100100111011101110111001101110001011101110111011000100000011101110001011101110111001101110111011101110100011101110110011101110111011000010101011101110111011101110010011101110110011101110111000101110111011101110111011101100110011100000111011001110101011001110111001100100111011000110100011101110001011101010111011001110111011101110111001100010110011101000111",
		"01100001011101110111011001110101010101110111011100010111000001110111001001100000011101110100011101010111011101110100011101110110001001110111010100010111011001110111011101010000010001110111010101000000011101100111011101010111000001110111010000010111010001110111010001110000001101110001011001110011001101110010011101110010011101110111011101110111011000010111011101110000011000110110010101110111001000110111011101100111011101110111011101000001011101000111011101110110011101110010001000010111011101010111001000110111",
		"01110111001101110101010101110010001001110000011101110100011100100001011001110001001101110100011101110000001001010111011100010111011101110000011101110111011101110111001000000111010000010111011100000111000000000010011101110111011101000111000001000011011101110111011101000001010001000111010101110111010001010111011101110111000101110111011100010111000001000111000100100111011101110111011101110011011101110001011101110000001000000111000001110100001000100100011101010111011101110110011100110000011101110100001001110111",
		"00010111000100100111011100100111010001110011000000000111011100100111010001110110011101100111010100100111001001110111011101110111011101110011011001110111010100010100011101110111001001110111011101110111011100100111011100010011011101110000011101110110011101110111001101110001011101110111010001110111001101110111011101100111000000110111011101110110011101110111011101110011011101110100011101110000011101110110001101110111011101110010010101110001011100000111001101110111011100010000011101000110011101110111011100100111",
		"00100111011101110111011001110111011100000111011101110110011100110111011101110101011101110111010101110111001001110111001101110100011101110111010001110111001101110111001101110100010101110101011101110111011100010001010001110010000000100111010101100111000001110111011001110001011101110111011101110111000001110001011101110110001001110111011101010111011100100101010101110011010100110111010101110111011100110111010001110111000001110111011100100111001101110111010101000111011101110111000001110010011101110011000001110111",
		"01100011000000000010011101010111011101110101011101110010010001110111010101110000010101110110011101110011011101110101000101000110011001110100010001110100011001110001011101110011011101110001011101100111011101110110011101100111001101110111011100100111011101110111010101110011010001110111010101110001010101110111011101100111011100010111001001100111011101110101011100100101011101000010010001110001011001110010011100110101001001100111000001110111000101100101001100010111000101110100011101110111011101110111011101110011",
		"00000111000101000111011100110010000101110011011101110111010000110111011101110111000001110101011101110111001000100101010101110000010100110111011101110111001101110000011001110100011100100011011000010010011101110111011100110101011101110010011101110111011100000111011101100111001101110101011101100011010001110110011101110111011001100111011101110111000001110111011101110100010101010111001001110000001000000111011101000001011101110111011101110100000001010000011101010111011101110111011101110001011101110101010101110101",
		"01110100010101110111000101110001010001110111011101110111011100000111011101110110011100110111011100110111011001010111010000000101011101100111010001100101011001110111011100110001000101000111011101110111010001000010011101110111011100110101011101110111011101110111011101110101011100100000011001110100011100000111001101110100001100100010000000000000011100000111001101110101011101100111011101110100011100110111010001110111011100100111011101110111001100100000011101110111010100000111011101010111011101110101000001110000",
		"01110111001101110100011001110111000001110111011100100001011101110001011101110111010101010110011101110111011101110010010001110100000001110001010001110111000101110110011101110111011101000111011101110111011101110010011101110111011101110001011100000001000001110111011001110011011101110111011101100111011101000111011101110100011100100111000001100111011101010111000000010111011101110111011101110101011100110111000101110111011101010000010101110111011101110010000001110111011101110111001001010000001000000111011001010111",
		"01100111000100100010011101110111000000000111001101110010010101110111011001110110011100100100011101010111011101110111011101110011011101110111011100110001010001110001000101110111011000100111001000000111010101000111011101110111000001110101011101110111001000100111011101110110000000110101011101110111011101100000011101110111011101110111011101110100000101110111011101100111011100100011000001110111011100000101000001110010000000000111011101110110010101110111011100100111001001110100011101110110011101110111011101110000",
		"01110111010101110001011101110111011101110101011101110111011100010111010100000111000001110100011100100111010001110011011101010110011000000010011101110110000001110111011001110111000101110111011100010110001100000001011101110111011101000111011101110011000101000111011101110111010101110111011101000011001101110111000100100111011100010111011101110111000100110111011100110111011101110111001101110001000001010011011001110111010101110111001001100110000101110111011101110111011101010001011100110111011101110101011101100111",
		"00110111011101110111001100010111010001010110000101110101011001010110001001110111011101010010011100110111011100100111011100010111011101110001011100000000011100110111000000100100011001000010010101110111010000000111000101110111011101110111011101110111011001110111011101110000010101110100010101110110011001110010010001110100011101010111011001100111001001110011001101110100011100100111011101110111011101110111011100010101010001000111011101110000001101110111011000110100011101010111011101110111011100110111001101010111",
		"01110111010101110111001000000010011001100000011101000000001101010101010101110100010101110111010001010001011101110110011100000111001101000111001001110111011101010111000001110111000001110111001101110111010001010111000101110111011101100111011101010111011100100111011101110111011001110111001101110111011101110100011101010111011101010111011101110111011101010111011101100100011001110111000001110001010001110111011101110000010000010011010100110111011101110111011101110111001100000011011101110111010101110111001001110111",
		"01000101011101110010010001000100000001110111000001110110010001110100011101110101010100010001001101110111010000110111001101110111011101110111011000000001011101110111011101010101011100010000011101110100010001110000011101110000011101110111001001110111000000110111011101110111011101110111001101110111011101110111001001010000011101110111011101110101000001100111011101110101001001110111011101110111001001110111011100110011000000110111011101110111010001110111011101110111001101110111011100010111011101110011011101100111",
		"01110001011101110000011101110111011100000110010101110011011100110111011101110111000101110000000101110111000101110111010101010001011001110111011101110111011101110111010001010111011101110111010001100111011101000111011101110111011100000101011101100111011100010111011100000111011001110001010001110111011101110110011101000110011101110100011100010111010101110100010000110011010001100000011101010110011001010111011100100110010001110111000101000111011100000111011101110111011100000110010101110011011101110111011100100000",
		"00100001011101110111011100100100001001110111001001110111010001110111001000100111010101100101001101110101011101110111010001110111011101110111011101110100011101000111010001110111010101110111001000010011011100110010011101110111011101110111011101110000000101110111000001010111011100110110011101110111010001100010011101110011000001110111011100010111011101110000011101110111010001010111011101010111001001110110000001110011011100110111000100100010011101110111011101010111001001110111011101110110010100100101011101010111",
		"01110111001101110111011101110101011100000110001001110111011000110011011101010111011101110100011101110111000100110111010101010110011100010111011101110111001101110111000100010100011100010111011101110011000100110011011100000100001100100111011001110101011101110111000001110111011101110111011101110111000101110111011101110111010000100111010101110101000001110110000100010111011100110100011101110111010001110001011101000111011100010101011001100111011101000111000001110111011101110000001101110011000000100001011101100100",
		"00110111001000000000011101000101010000110111010001010110010001110111011001000111001101000100011101110111011101010111000000110111000000010001011101110111011101110001011101100101011101110001011100110011011101100011011101110111011101100111011101000111010101110111001001110001000001110111011101000110000101110111011101110111011101110110001001110111011101000111011101110111011101000011000001110111011101110111011101110100000001110111010001010101000101110111011101110010011101110001000101110111011101000001011101110111",
		"01110111001101010111011000010101010000100110011000110011011101010011011101110100011101110111011101110111000000000111011101110111010001110111011101110000000101100111010101000001011000000000011101110000011100010000011100110111011100100011011101110111011101110111011100100101000001110111001001110111011100110111000001110111011000100111000001110111010001100111010001010111011101100111011101110101011100010010011001010001010001110111010101110111011101110101011001110111011100000111011101110011011101110111011001100111",
		"00100111011101110000001001110111011101110111011101110111011100110111001001110111011101110111010101110111000101110111010001110011001101110111011101110010011101110111010001110111010101110111011101110010000001110111000101110111000001110110010001000000011101110100010001100010011101110111010101110011011101000010000100010011011101110111010000100111011001110111000001110111011101110100011101110100001001110111011101110010011001110011010000110111011100010111011101110000011100010111000001110111011100100111010101110110",
		"01110100011000100111011101100111011001100000011101100000011101010111000001000111011101100011010001100111010101000111011101110111011100100011011001110111011001110011010101110110001101110111000101110111000101110110011101000111001101110111000100000111000001010111011101110000011101110100010101100111011101110110011001110011011100100111011101110110011101110111011101000011011101110111001101110110011101110111011100110100011101110101011100110000000100000000011001110001011100110111011100100111001001110111011101110101",
		"01110111000001110011001100010111011101110111011101100111011101000000011101000111001001000011011100110000001100110101010101000110010001010000010001110100011101110111001001110000000101110001001101110111011101110111011000110111011101110110001101110110011101110011001001110001011101000111011101110110010101100101001000100100011101100001011001110110011101010111011101100111011101110111010001110001001001100111011101110011011101010011011101100010011001110111011101010111011101110111001001110101011101110111000001000011",
		"01110011010000010111001101110111010100000011001001000010000101110111001000100111011100010110011101110010011101010111001101110111011100010111011001110111011101100000000101110110011101110111011100100011011101110101011101110000011101110101011101110010010001110111000101110111011001110101010101110100011101110110011100110111011101110001010101110111011001110001011101100111000001110000011100010111011101100111011101110001000001110101011100000011011100100111011100110111000001110111011101110010000100110111010100110111",
		"00100111000001110111011101010110011101110111010101110111001101100111011100010110010001000111011101110100011101110111011100110010011100000001011101110100001000100111011101110111011100000111011101110111001100110111011101100111011101110010001101110100011101100111001101110111011101110111011101110011011101010111001001110101011101110111011101000111011100000000000001110111011101110101011100110111011101110111010101110111011101110111000101110111011101110111001000000111011101110111011101110111011100110100011101110101",
		"01100111011101000111011101110111011101110111011100000111010001000001011100010101010001100111010101110111011101110111010001110100010001110111011100110111011001110010011101010111011001110100011101110111011101110011000001010010011101110111011101110111001101110100001101110010011001110011011101110111011101110000010100010010001000110111000001110111001001110111011101110111011101110111000101110000011001000101000101110101001101110111011101110001011101110111000001010111011101000111001101110111011101100001011101010111",
		"01110011011101110101001000000110010101110111011101110110001001110111011101100100011101110111010001110001011101100111010101110010011101110111001001110111011100010101011101110111011101110111011101110111011001010001001100110111010100110111010001010111011101110010010101110111001100110111010100100111011100100100011001110010000001110000011101110111010001110111011100000011010101110101011101110111011101010111001101110111011101100111011101110111011101000001001001110111011101110101011100110011011101000111011101110111",
		"01110000011100100010001101110000010101110011010000100100011101110000000001110111011101000111011101100001011000010111011100100111000001110001011101110100011101110111011101110111011101110111011001110000001101110111011000110111010001110110001100100111011101010001011101110001000001110110010101110111010000010101011101000111011101110111010001010111010101100101011101110011011101110001011100100111011100000011001101110100011001010010011001110010011101110000010101110100011101110111000000110000011101110111011101110111",
		"00100110011101110111011100000111011101010111011101000111010001000001001001010000000001110111000001010010010101110100000001110000011101110111010000000111010101000111000000010000011101010111011100100001011101110101011101110111011101110111011101110000011100000111011100110101010001110111000001110010000000010010011101110001011101110111011100110110010100110111011101100111011100110000001100000011001100100111010001110011011101110000000000010011011101010011011101110101011001110111000100000111001101110111010001110111",
		"01110110011101010111011101110111010101100111001001000111011100010101011101110111011101000111011100000100001001110100011101000111011101110111011101110100000101010111011101100110001101110111011101010111011101010101011101110111011101110111011100100111011100110111011101010111011100100111011100010010001101110100011101110110010101000101011101010011011101100010011100000000001001110111011100000100010101110111001001110111001100010111010101110111010101110111001001110101011101110100011100100001001001110111001101000110",
		"01100110011101010110011101110101000001010111011101110111011101110111011101110101011101110111011101110000011101110111011101110100001001110111011100100000001000010010011100110111011101000111011100100111000101100111011101110111011101000111011001110101000001110100011101110011011101010111011101110101011101010000001001000111011100100001000000010110001101110101000101110111010101110001011101110111011101110110011101110111000101110111011100110111010101110111011101110111011000010111011101110111011100100000010001110000",
		"01110111011000100101000101000111011101110100011100010111010100110111011001000110011101110010011100110010011101100111011101110010011101010111001001110111001001110111000001110100000101110001011101110101000101110111010101100111011100100111011101110101010001110111011101110000011101100111011101110001000101110001011101110100001100010100011101110010001100010011011101110111001001100101011101010111011100110111011101110111011101110111011101110111001001010110000101010111011101100010011101110001011101110111011101110111",
		"01110111010100010111011100110101011101100010011101110111011100010011011101010111010101110111000101110111001001110010000101110101011100110111011101010100011100000111011101110101001000010111011101010011011101110011011101110111010101110111001101110000010101110111001000000111011101110111000101110100011101110001010101110111011100010001011100100100011101110111011100000001001101110111000101010011011101110111000101110111011101110111001101110000000001110111001001010111011001110111011101000000001001010111011100000000",
		"01110100010001110010011100010101011101110101011100000111011101110111000100000111001100100111011101110110011100100101011000110100001101000111011001110111001001110111011101110111000101110001011101110111011101110111010101010111011101010111000001110000011101110010010001110010010001110111001101110001011100110111011101000111011101110010001100010111001100100001010000110010011101110111011101110001011101110111011001110111010101010111000001110001010001100001010101110011011101110111011101110111011101000110011100000111",
		"01110111011100100111010101010100011101010111011101110011011101110111010001110111001101010111010001110010011100010011011101110111011100000010000001110111011101110111011101110111011101110111000100110111011101110001011100110111010001110111011100110110011101110100011000010000000100010111000101110100010001010111011100000011001001110100000100110111010001110111011101110011011101110001010001110111001101110111011000010011011101000011011100110010011101110111000000000111011100100111011100110000011101110111011100010100",
		"01110011000001010000010000100011000001100111001001110001010100010111000001110111011101010011011101110111011101110001000001110111011101010111001000010011011101110111010001110111010001110010010001110111010101010111001100000111000100010111011101110011011101110111011101110111010100110111011101110111011100000010001001110111011101010011011100010111011101100101011101110110011101110111011100100111001001110111011101110111011101100000011100010111011100000111000001110111000101110000011101110101011101110110010000110011",
		"01110010011101110101011101110111011101110001010001100111000000100011000100110100011101100111011000010111011101100111010100000111011101000111011101110111010100010111011101110111011101110111011101110111011101100111001001110000011100100010011001110111000101010111011101110111011100100001000100110101001000110011001101110111011101110101011101110111011100000111011001110111001101110000011101110110010101110111011101100111011000000111001101110011001100010110011101110110011101110111011101000100011100000001011101110001",
		"00100001011101110111011001110111000101110100011100010011001001110111000100010111000001110000011101000110010100100111011101000100011101110111010001110001000101110001011101110111011101110111011100000110011101100000000001110110011001110111011101110111011101110100010001110111010101110111011101110010000001110000001101010000011101110000011101110111011101110001001101110111000001110111011101100111001001100111011001110110011101000111001001110111001100010111010001000111010100010111011100000111001101110001011101000111",
		"00010111001101110100011100100010011100100111010101110111011101100010001101110110001101000110000001110111011101110111000000110111000000100111011001110110010001110110011101110111011101110111011101110101011101110111011101110111001101000010011100100111001000110110011101100111011001110100010001100111011100100111010001110000011101100000000101110111010001110111011101110000011101100111010100000101010001110111011101110101000001110000011101110111011100110101000100000010011101000010011100100110011101110001011100010111",
		"01110110011101110111011101110111011101110111011101110100011100010000011100100111011101000111001101000111011101110101011101110000001100100100011101000111011101110110011101000000001100000111010101110111011101100011000001110011010001000111001101110111010001110111011100100011011101110111011100100111000001110111011101110010011100110111011101110111010101110111010000110111010101110111011101110111011100000111010100110111011100010011011101000000001101110001010101110111010001100100011101110011011101110111011101010111",
		"01110111011101110111011101110001011101110001010001110111000001110010011100000111011101110010001001100111011101110100001100110100011100000111011101110000001001010111011100010111011100100111011101000111011101110111010100110001011001110000011101110010001101110001011101010111010000100111011100010010011101110010000101100111011101000111010001110111011101110100011001110111011101110010001101000111011101000111011100110111011101110111011101110110011101110000010100000010011100100001010101110111011100000110011101010111",
		"00100110011101110111011101100000011101110111011001110101010001110111011100000010001101110111011101000111011101110111001001110111001001110111011001110111011100010111000100100111011101000111011101110010011101010001010000010111001101110111001000010001011101110111010001110000011101110111011101110111000101110101011101110111011100110111011100100101001101110010010101110101011001110001011101110100011101110111011101010111000101110111001001100111011101110111010001100111010001000000001101000111000001110111011100010111",
		"01010111011101010100011101010001001001110111011101110001001000000111010101110111000101110111001101110010011101110111011101010111000101110001011101110101011101100100000101000111001001110111011100000111011001110001011101110011001001110111011101110011001101110001001000110111000001110111011100100011010001110111001101110111010100010111011101110111011101000001010001110111000101110011011101110111001000010111001001010100000100000111001101110010011101110111011101110010011100100100011100100111011101110000010100100001",
		"00010111011101110111011101110111001101110111011101110111011101010111000101100100010001010001011101100111011100010111001101110111010000110111011100100111011101110001011101110111001101110011011101000111011101110011011000100111000101110111011100010001011100100111011100000111010001110101011101110011011101110000011100110111011100000111000101010111011100110010011101110111011101110111000100000001011101110111001101000111011100110111011100010111010000010111001101110111011101100111011101110111001101110111001001110100",
		"01110100010101110111011100100011011100110111001101110000011101110111011101110100001001110111011101110101010100000111010101110111011100100111010001110000011101110001011100110111010100000111011101110111011101110110001000110101011101110110011101110010001001110110010001110110011101110111011101110111011100000011011101000111011000100110001101100111011101110111011101110001011101110011010000000111010001110111011101110111011101110001011101000111011101110111011100010011011100010111011101110000011101110111011100110111",
		"01110111000001110111011101110111011101100111010001000100011101110100011101000011011101110111011101110111011101110111011001110111011101110100011101010101000001110111011101110111011101110111011101010111011101110111000101100111001000100101000000010111001001010001011101000111000100010110001100100111011101110010011101110011011100000010001100100000000101110111011101110110011100110000000100110111010000100111011101110101011101110001011100100100010001110100011100000111011101110000010101100001010101110111011101110010",
		"00000111000000100111011101110001011100100000011001110111000100000111000001110000011100000111011101110111010001110001011101000111011101110111001001110111011101000000011101100111011001100111011101100010011100100000011101110111010000100111011100110001011101110100011100010110001000000111001101110001011100000101011001000111001001110111011101010111001101110111011101110100000000100010001101100111011100100111011101110111001101110111001101110111000100010111011101110111011101110111011101110111011101110111011101110111",
		"01110111011101110011000101100010010001110111000100000110000000000111000000100000011001110111011101110111001001110111011100110100001101000100011101100000001101110010010001110111001101110001011100010111011101100111011100000101001101010111011101000111011100010111011101110111011100110111001001100001010001010111011101110100011100100111011100110110011101110111011101000111000001000100011100110111001001110111011001010111011101110111000101110111010001110001011101110010011100100100011101110101011000010100001101110111",
		"00000111011101110000001001110110010100100111011101110111000100010101001001110111011101110111011000110110000001110111011100110111011101110011010001110111011100010111011101110111001001110010011001110101011100000111011101010100011101100111010101110111011001100000011101110011011101110101011101110111000001110111011101110111011001110101011101110111010001110111011100110111011101110111010001110010010001000101000001010110011101110010000100010100011101110010010001110101011100000110011101110100011101110000011100000111",
		"00100010011100110101011101110111011001110111011100000111000001000000010001100100011001110100001001110111011101110111011101110111011101110111000101010010011101100101001001110111011101100111011101110010000101110000011101110000000001110100001001110001001101110001010101110111011101110010011101110100010100110111011101010000011101110011001101110011011100110111001001110111010001110111010101110011011101110111011100000111011100110111011101000111011101000000011101010111011101000111000101110100011100100110001001110111",
		"01110111001100110111011100110111011101110000011101110111000100100101011101110111010000000010011100100000011101000110011101110111010100100111011100100111011100110011011101110111001100100111011101110010010000000111011101110111011100100100011101000100011101110111011100000001011100010111011101110111011101110100011101110111001100010011011101110011001101110111001001110111011100110011011101110101011100010000011101110111011101110111011101110111011101110100000001000111011101110111011100000111011101110001011100000111",
		"01100111011100100011010100010111001101110010001001110001010101110111011101110111011101010001011100010111001101110111010001010111000001110111011101110111011101110110011101110111010001110111011101110101011001110100011101000001011101110111011101110111001001110111011101110000011101110000011101100011000100000111000001010111010001110010011001110011000101100011000001110010011101100011010001100101011100100111010101100111011101110111011101110111011101110111011101110000011101010111010001110111011101000111000100000000",
		"01110111011100000100011101110111000101010010011101110111001001110111000101100111011101110111011100100111011100000111001101110011011001110111011101100100010001110111010100100111000100010111011100000111011101110111011101110111010001000010011101110001011100000111000101110111011101110100001001110111001000100111011101110101001100000111011100010111011101110111010001110100011101000001011101100111001101110101011101110111011001110111011101110111000101110111011100110111011101110111000001000011011001100110011101110111",
		"00000110000101110111010000100100011101110001011101110111011001110101011101010100001101110111011101110011010000110111011001110111011101110001000101110111011101110111000100110111011101100111010000010001001000110111000001010111011101110101011101110100010101110001011100110111011101110111011101110011011101100111000101110100011101000111011101010111011000010111000001110111011101110110011101110000011101110100011101110110011101000111001101100111000000110111011101110010011101110111010101110111011100000011011101110111",
		"01110101010100000111011100000111011101110000011101110111011100000111010101110111000000000111011101110000011101110111011101110100011100010100000101110000011101110101000101110101011100110111011101100110011100100010001001110010010101110111011101010010011101110111011100110111011100100111011100100111000101110111011100110111011101110111000001110011011100000111011100110111011101110111000001100111011101110111011101110100011101000001011101010110011101110111001101110010001001100111011101000111001101110011011101110111",
		"01110111011100110111011101010111001101000001000100010111011101110111001001110111011101100111011100110001011101110011001001110110000101110111011101110000011101110111001101110010011101110111011101110100011101110111001000000001010001110111011101110111010101110111000000110100010101110111010100100101011100110111010001110010010100100010011101110111000001110111011101110111011101110111011100000100011100000111000001110111011101110111010001110101011100110111011101110111010001110111011101110111010001110111011101110111",
		"01000111011101110111011101100001010001110111011001110110011100010011011100000011011101110110011101110010011101000111011001110011010001110011001000000001011101010011011101000111011100010111001101110111011101100001011100100010011100000101011100000111010001110111000001110000010101110110001001110111011100100100011101110011011100100100011101110001011101110111001001010100011001110101001001110111011101110111011101110111000101110111010001110111011101110111011100010011011101110111011101110111011101110011011101110101",
		"00110111011101110100011101110111011101000100000001110111011101110000001001110111011101110101011101110111011100110111011101110001011101110111011101010111011000010111011101110110011101110111000101110110010001110100010001000011011101110101011100000010011101110111011001010010011101110011010001110111001000110111011101110111001001110111010101100111011001110010011101110110011101110111001101110111011100010111010001110001011100000001000101110111011101110111011101110111011101110000000001000010011101110111011101110111",
		"01110110010100100010010000100111011101110010001100100011011101110111011101110111011101100001000001110111011001110111011101110010011100010001001001110111000101110111011101110111011101100000010100010111011000100111001101110111000001010010011101010111010001110100011100110111011101110011011001110110000100100111010001110100011100100010010100000111001001110111011101110111011101110111000101110010011101110111011100000111001001110000011100100111001001110110011100110111011101110110010101010111011100110111011101110111",
		"01110010000101110111000001110111000101110111011001010111011100000001000001110100011101000111011101110111011100010111011100100111001101110111011101100001011101110101000101110101011000110100011001110111011101000111000101010111011101000111011100000101011001110100001100010111000101110111011100000111000001100111011101110111011101110110000001110111011100010111011001110111010101110111000001010011011101110111011101010000011101110111011100100111011101110011011101110111011101110101011101110111010001110111000001110111",
		"01110110011101000111011100110010011101110111011100100011011001010111001100000111011100110111000001110010010101110010010001100111011001110100011101110010001001110011011101000111011101000111010001110010011101110100011100010001011001110011011101110010011101110110001001110001011001110111011100100111010001110111011100010111011101110111011101110110000101110111011101110010011100010110011101010111010001000111001101110111011100100111001000100101011101110100011101110111011100000111000101010101011101110011000100100110",
		"01110101011101110011011101110111011101110010011001000111010101110111011101110111011101110011010001000111011101110111011100100111011101110011011101110000010001110111011101110110011101110001011100100111001101110111011101100111001101110111011001110100011100010110000001110100011101110111001001110111011101110111011100100011011101110111001101110111001001110111011101110111011101110111011100010100011101110111011101110111010100000111011101110111010101110111011001110000000001110100011101110011010101110011011101100000",
		"01100111011101000111011100100110000001100111010001110111011101110111000001100111000101110100011001110111011101110010001100000010011101110111000101110111010001110101011001110111001001110111011000110111011100100101000101110110011101110111011101000011011101010111011101110111011101110101011100000111011100110111011101110111011101110101011101110111011101110111011101000111010001110111011101110111011100110111011101110110000001100111011100010111011101110101001001110001011101110111000101010010011001100000011101110111",
		"01110111011101010111000101110001011000110111011100100111000101110111010001100111011100000100011001110110011101110010011100100000011101010111011001110111011100110001011101010111011101110111011100110101011101110111011101110111001000110010011101010111001001110010000001110111001000110101011101110111011101110111011100110001011101110101000101110010011101110111001101110110000001110111011101000111000001110111011001110101011101100010011101110111001001110111001101000101011101110111000101110000001100010110010001110001",
		"01110011001000110101011101110010011101110011011001100101001100100111011101110111011101110111011101110111011101110111010001110111001101110110011101010111011100100110000001000111010101110101011001110010010100100111011101110111000001110110000101110001011101110111011100100111010101010111011100100101011101110111011101100111011101110111011101110111011100110111001101110111011101110111011101110101011100010111011001100111011101110111011101110111011100100111011100100111011100110111010001110111001001110111011001100111",
		"01110111001100110100000000000101001001100111011101110110011101110111011101110111011100100010011101110001011101110011001100010111011101110010000101000111011101000111011001010111011101110111010101010110001100000111011100000000011101110111001001110111011100100010011100100111011100000111011100000100011101110111001100010111011101110101011101110111011100100111011001110111010101110111011101110111011100100111001101110011011101110111011101010111000101100110011101100001011100110100001001110111011101000111001000110111",
		"00010110011100100111011101110011001100100111011101110011010100100011011101110110011100000111001101110010001101110111011100000111011101110110011001000111011100000101011001110111011100100111011000010111011101110111011101000111011100010111011101110111011101110011010101110011011101100111011100010010011000110111011101000110011101110111001001110111011101100111011100100000011101000111000001010111001001010111001100000010011101100111011100000111011101000111001100000111001000000011001100100111011101110101011100010110",
		"00100111011101110010010100110111011101000111011100000111011101000111011101110101011101110101011101110101001101000101010001110111011101110111011100000111010101110111011101110111010101010111010000100111011101110000000101110111010101110111010000010111011100010111011101100100010001110111011100110011011101110010010000000111011100010111011101110100010001110010011100100111011101110101010101110010011101110110011101010001011100010111011101110110011101110111011101110110011101110000011101110110011101110101011101110010",
		"01110111010101110111011101110000011101110111011100100000011101110111000101100100000000000111000001000111011101110111011101110111011101000111000101110111011101110010000000100111011101110101011101010100011101110111000000100111000001110110010100110111010101110011011100010110011101110111011101110111011101110111011001110111011001110111000001110111001101110000011101100111011101110111011101110111011101110100000101110111000100100001011101100000011101100111011101000111001100000111011101000111011100110111010101110010",
		"00100111000001110111011101110111011001000111011101110111011100000001011101110010011001010010000100100111011100010111011101110111011101110111011101110000001001110100011101110011011100100111011101110100011001110111000001110111011100010000010001110010011100010111011101110111001001000001011101110101011101010111011101110110011101110111001001110111011101110111011100100111000101110100011100000111000001110111011100010111001101110111001000010111011101110111001100110111011101110111010101110111001000100100011101110000",
		"01110110011100110111011100000111011101110111001001110101011101110110001001110111000001110111011101000110011101110111011101110100011100000100011101110001011101100111011101110010011000010011011101110111011101110011011100010111011101100101011101110111011100010111011100010111011101110111001001110111010000100011001001110111010001110111001000010010011101110111010001100111011101110111000001110111000101110000011101000111011101110001011101000111011101110111011101110111011101110111011101000111011101100111011101110000",
		"01110110011100110111011100010111011101110111011101110111000101110110011101110111000100110111000101110111011101110000011100000111011101110111010001110111001101110110010101110111011101110111010101100111011100100111000000010100010100000011000001110011001000010010011101100010011100110111011001110010001001110001011101110111011100000111011101110010011100100010011101110100011101110111011101110111011101110111011101110010011001110111011100010011010000110001011101110100011101110111011101110111011001100111000101110101",
		"01110111011100000111011100010000010100100111010101110000011101110111011100000001011001110111010000110111011001110111011101000110010001110111000100010001001101110111011001110111011100000000011101110111010101110111011101010001000001110111000101110000010101100111011101100111011101010001011000110111001001000111001001110111011101110111011101110101011100110010011101110111000101110111011101110111011101110111011001110111011101110101011101000110001001110101011100110010010101110110011000110111000001110001001000110001",
		"01110111011101110100000101000100001001110111011101110111011101110111011101110111011101110111011001110111010001110111001001110000011101110010010101110111011101110001011001110101011101110011010001110111011101110001000100110101011101110111000100000111000000110101011100100110011101110111011100000011011101110111011101110110011001110111001001110111011101010111010001110010001001110110011101110100000001000111011101110010010000000111011101010111011101110111001101110111001101110101011101110100011101110101011101110000",
		"01110111011001110111011101110111010101110111011101110110001000110111000001110011011101110111000101110011011000000111000100100000001101110111011101100010010001110111011000000101011101110101011100010111011101110111011100100111011100100111011101110111011101110100011101110000011101110111000001100111010101110111011101100101000001110110011101110111011001000111011101110110010101110011011101110100011101110010011101110111011101000111011101110111000101110100011101110000011100010011011101110100011101110111011101000111",
		"01110111011101110111011100100100011101010100011101110111011101100111011001000111011101110111011100110110011101110101011100010000011100010010000001100111011001010011011100010111000101110001011101110111010101110001011101110111011101110111011101110111011101010111011100010111011101110110010101110011000100110100011101010111011101110100011100000111010000110111011101110111011100100000011101110111010101110111011101110111010101110111011001110111000101110111011100100111011001110111011101110110000000110111011100000100",
		"01110000011101110111011101110111011001110111011101110101011101110111011101110001000100000011011101100011011101110011011100110111001101110111010101110111011101110111011101000111011101110111010101110010010000000011010100010101011101110011010000100111011101110111011101110111001101110011011101110100011101110100011100000111011100110100000101110001011101110010011101100100011101110101000100110100011101110011011101110100010101110111011101100111011001110100011101110111010001010111011100000111011101110010011101110111",
		"01110110011101000111001001110100011101110100010000100101000001110011011101110010010101110111000100100111011101110111011101110001011100010010011101000011011101110111011101110111011100010101011101110111011101110110001000100111000100110001011101110100011100100100011101110111011101110100000101000111000101110111011101110111011101110111010101100110010001110111011101110010001100110111011100100000001100000110011100000010001001110011011100000111000101110011000001110010011100110001011100110111011101110111010001110110",
		"01110111010100010111001101010111000001110111001101110100011101010111011101110100011001110111010101010111011101100001011101110111011101110000011100110001010101110111011101110100010101000111011101110111000100100111011101110111011101110111011101110111010101110111000101110111001001010101011101110111000000010101011001010010011101110111011101110111001001110111010001110011011001110111011101110111011100000110001101110011011101110111011100110100011101110000011101110111000001110000011101110111011100110011011101110111",
		"01110111011100010111011101110111011101110111010101110111001000010110001101110100011001110111011101110111011100000100011101110111011101110111010101110111001000010110011101110011000101110111001001110111011101110111010101110011011100000101011101100111011101110010011000000111000001110110011101110111011100110111011001110111011101100011011101110011000101110111001001000111011101000111011101110001000101110111011101110111000101000111001100100111010101110111011101010111011101110110011101010101011101110100011101110111",
		"01110001011000010111011101100111011000100111011101110111011100110111011100010111011100100111011100000110001100000111010100010111011101110111011100110111011101010000011100110110011101010010011001100111010001000100000101110111011101110111011101010101001101110001001001110111000101110010011101110110011101110111011101110000000001110010011101110010011101110111010101010111011101110111011101110001011101110101011001110110001101100111011101110111011100010111011101110111011001110111010101110111010001110111011101110111",
		"00110000011101110111001101000111010001110010011101100011000101110111001101110111011001110111001000100011010101110011011100000111011101110111001101100100000101110110000101110110011101110111011100000101011101010000010001010111010000010111011101010111011101110111011101010111001101110001010101000111011001110111001001110111011101000111000101110111011101110111011101110111001101100111000001110111011101110111010101110111011101100011011101110111011101010110011101110010001001000111011101110001010101110111001001110111",
		"00110010011101010111001101110110011100100111010001110111001001110100011100110101011101110111011101110111010100000110011101110111011101110111011101110111011101110111011100000101011100110111010000010111011101110111010000100010011101110001011000110101011101110111011101110110001101110111011101110111001101110010011100110110011100100111001001110100001001110010011101110111011001100010001001110111011101110111000101110011011101110111011101110100011000010111011001110111011100010000011101110111011101110101000101110111",
		"01110111001101110111011101110111011101010111000101110110010101110101000001110111011101110111001001110100001101110111011101010111011101000000011101110111011101110111011101000111011100010100011101110111010001110111011101010011011101110101011001010111011101110000011101110010011101110111001001110101011101110001011101110111011101000111011101110011011101110111011101000111011101110111011101110011011101110111001101000111010100110000011101110111011100100111011100110010011001110111011101110111011101110011010101110111",
		"01110111011101110010001101110111011100100010001001110111011100110010000101110001011101110111011100100111001100010111011101110111011000000000011101110110011101110101011101110011011101100110011101110010011101110011011101110111000101110111010001000100011101000111001100000111011101110111001100000111001000100111011101100111011100100111010001110111000101010111010101110111000101110111000001110000011101110111011101110111011101110111011101110111011101110111011101110111011101110000011101100111001000010111000101100111",
		"01110111011101110010000101110000000101110111001001110000001100110010011101110111000101110111011100010111011101110111011101110010011101010101011101000111011001110111011101110110010000000111011101110111011101110110011100110001011101110111011101110111011101110111011101010100011101110100000000100111000001110111011101110110011101110010011100100111010100110000000101110011011101110111011000110111011101110111000101010101001001110001011101110110011101110111011001010001011101110111011101110010000001110111001100100110",
		"00010101001001110110011101110100011101110001011100110111011100010111000000100011001001110111011101110111011101010111011101110000011100100101011001110111011101110111010100000111011101110111011101110111011100000111011101110011011101110100000101110000011100110100011101110100011101100100011101110111011101110001011101110111010101110111001101010111011101110111011001010111011000010111011101100111011101110010011100010011011101110001011101000111011101110111000001000101000101110111010001100011001001110100000001110000",
		"01010111011101110001011101110010011100100111010100110111001101110011011101110111001001110001001100000101011101000111001101110001011100110110001001110111011100010111011101100010011101110111001001110001011100110001011101110111011101000111011100100000011101110111000000000111011100010111010100110010011100010001000001110111001001110111000000100111011100110100011101110111000001110111011101110111011101110111011101110101011101010111001101110010011100000111000000100111011101110111011101110011010101110100010001110111",
		"01110111001001010111011101110110000101110111011101110010011101110001011101110111011101100111000001110000011101110111011100000111011100010111011101110111000001110100000001110100011101010111011000010111011101110111011101110110010001000111011001110111010100010111010100110111000001110001001001110111001101110001010000000100011101110001001101110111011001110111001101110000001001110111011001110111001101110111000001110101011100000011011100110000011101110111011100000111011100000101011101110001011101110111010101000111",
		"01110010011000010010000001110111011101110111011000010000011100110111011100010110011101110111011101110111000100110111010000010111011101110010010001000111011001110110011100100111001100100111000101110111011101110111011101110111011101010111011100100110011100000011011101010111001001100111010101110111011101110110000001000010011101110110011101000111001001110011011101110001011101000111001100000111010000010111011101110011011101110111010101010111011101010111011101110010011101110111001101010111011000100111011101110010",
		"00010101011001010111011001110001011101110110011101100111000101110111011101110000001000000111000101110111010101110011001001110101000100010111001001110111011101110111010101110111011101110011011100010111000001100111001000100001010100100000011101100000011100110111000101110111011101110110011101110111010001110111000001110001011101000111011101000111011101110011010101110111000101110111011101100111011101110001000100110010011101110111011101100001010101010101000000100111011101110011011001110011010101010111000001110011",
		"01110000011100000001011101000101011101110111011101000111011100010010010000110111011101010011010001110111011101110110000001110111011100000011011001110111011100110011011101110101011100000111011101110111011101110011011100010111011101110111011101110100011100100110011001110000001001110111001101010111011000100111001101000111011000110101011101110111011100110000011101100111000001110111000101110111000001110111011101110111011101110001011101000010011101110111011101110111011101110111011100010111010101110111001000000111",
		"01110011011100100111011101000111000001000111011101110110011101110000011101110110001101110111011100110101011101110010011101100111011101110111011101100111011100010010011101110110001101110111011101110001011101110000001101110111011101110111011100010101000100010001010101110001000101110111000000010111011101110111011100010100000000010111001101110000010101110100011100100101011101110110011101000111011101110110011100000111011101110111010001100111010101110101011101110101011101110110001100010111001001010111011101110011",
		"00010111011100010111010101110110000000110111011101010111010001010000011100110110001001010100011001110001011101110101011100100111010101110111010001000010001001110110000000110110001101110100001001110111010001110111010001110111011101110111011100110111001100010111011101100001010001000111001000000111011000100001011100110111011100100111001101110011011101110101011100110111011001110111011101110110011101110001010000010000001001110111010100100111001101110111001100110010011001110111001001110110011101110101011100000111",
		"01100011000001110111001100110011001101000111010001010111011101010111011000100011011101110111011101100111011001010111010001110101011100110000011000100101000001110111011101010000000001110111011100000010011101010111011101110111010000010111001000010111011101010111010001110111010101010111011101010111011101010110000000000111011100010111011101110001010000000111011101110011011100000111000101010111001001110111011101110011011101110110011101110001000100010111010001110111011101110011011001110100001101000111011101110110",
		"01110111011101110111000101110111011101110111011100110111000000010100001001110100011001110111011101110111011101110111010001110111001001110101011101110111011101100110010001110111011101110010011101110111011101110111011101110000011101110000011101110111011101100110011101110100011101110110011101110110011001110001011101110111001100010010010001110010011101110101011101110111011101110111011100100111011100100111011101110111001000010111001001110111011101000110000101110111011101110111011101110111001000100111010101110111",
		"01000000011100110010010000000111011001110111011100110111010001110000011000100110001101110011011101110000011100000011001001110111011101110111011101100111011101010011011100100111011100000100011001110010011101000111000000010111011101000010011001100110011100010000000001110001010101110001011101010110011100110011011101110001011101110110011100010011011101110111001001110001011100000111011101110111011100000111001001100111011101010101001000100100001101110000011101110111011101110111011101110111000001110010000001110111",
		"00100101011101110100010101110100001000100111000001110111011101110110011101010010011000100011011101100111000101110111010101110110011101110111001000110111011100010111000100110011000101110111010001110011011101110111011101110011000101000111011101000111010100100111011001110111010101110011001101110111011101100010011100000000010100100001001001110010011100100110001101110111000101110110010101110010010001110110011101110100001001110111000001010111011101110010011101100011000001110111010001110111011101110001000000010111",
		"01010111011101110111011101110101000001000111000101100111000101100111011100100111010101110111000100110101000001100101011100110101011100100100010001110111010001000010000100010111001001010111011101110111011101110110011101110111011100110110011101110111011101010111010001000110001001110111011101110111000101100111010000100011011101110111011101110101011101100010000001100111000100110111001000010111011101100111011101110111011100110111011101010000011100100111011001110111011101110001011101110000001001110010011101110001",
		"00010000000101110111011101000111011101010110001101110111011101110111011101110000011100000100011101110011011101110000000100010100011101010111011100100111010101000110011101110111011100000111001100100111010100000011011101110110011101100010011101110111011101110101000001110111011001110111011100110111001001110111011100100111011100010111011100000111011101110000011101000001011101110111011101110111011100100010011001110100011000100111011101110111010000000111000001110000011101100111001101110111011100110111000101000111",
		"00110111011101110111010001110100000000000111000101100111010101110111011101110111011101110010011101110011011101110000011100010011011100110101001101000111011100010111011101110111010101000110011001110110001100110000011100010011011100010110011101110111011000010110011101110111000100110001011101110111011100000101011101110111011101110111001100100010011101110111011101010111011101110010011001110111000001110111001101110010010001110000011101110010011101110111010001110111011001010110000001110111000101110001010101110111",
		"01110111000001110001011001110101011101110011011100110111011100100000011101110111011101110111000001110111011100110110001001010111011101110111000100110111011101000111001001000011000001100111011101110111011101110111001000110111011101110101011101100111001000010001011100000111011100100111011101110111011101110001011101110111010001110010011101110111001101110111001101110111011101110111000000010111011101110111011101010111011100010110000100000100000000110111011101100000011101100111011101110111001001110000011101110111",
		"01110111010001110111011101110110011001110001011100110111011101110010011101010010001101110001011101110011011101110111001001110101010000000101011101110011011100010111011001110001011101100011000101110010001101110011000101000111000001110101010101110011011101110111000101110111011100100111011101010011001101110011001100010000000101110110010000100111010101010111010001110000011101110111011101110000010101110111011101100001001101110001011100000111011101010110011101110100011101110111011100100111011101110010011101110101",
		"01110111001000000111011101110111011100000001011001110111001101110111011100000000011101110111011101110111001101110111011101110010011100000111011101110111011101000111011101110111011101000111011101110111010001110010011100100111010100000111000001110110000101000101011100010111011101110111011101110001000001110101011101000010011100010110011101110111011101110000001101110101011101010111001001110111011100100111011101110011011101110110010001110000001001010111000001110011010100010011011101110101001000110111010101000111",
		"01110100011100000111011101110011001000010111011100110110011000010111011101110111011101110111011100110100011101110100011101110000001001010001001001000001010101000010011101110111011101110111011101110101011001110111011100000111011100000010011101110111011001010111011101110111011101110111011101110111001001110111010101010000001000010001000001100111011101110111011100110000001001100100011101110001011101000011000101100101011001110111011100000111011101110111010001110111000000100111000101100111001001110111010100010011",
		"01110000011100100111001101110110011101110011011101110000011100100111011100000010011101110010011101110001000001110101011101110010001001110111011101110010011101110111011100100111011101110111011101110111011101110111011101110111011100100111000001010100011101110111011101010001001000010010010101110111011101110111011101110111010001110111011100010111010101110001011101110111011100010111011101000001011101110111001001000100011100000010011101110111011100010011011101110001011100100100011101100011011100110111001100100101",
		"01110111011100010110011100110100011000110100011101110011010100100111011101110001010001110111011101110010010101110111011101110111011101110111011001110111011101110001011101100111011100100110000100000111011101110111000001010111011101110111011100000010011101010111011101110111000000010111011100010000010001000111011001000111011101110000011101100111001101110111011101000111011101110111011101110100000001110001011101110111001100010001011101010010011100110111000000100100011100010100011100100111011101110111011100010000",
		"01110111011101110111011101110111000001000110011101000111011101010111011101110010011101110111001101000111011100010111011100010101011101110111011101110010000100100111011101110111011101010111011101110110011101110111000001110101011101110111001001110111010100010111011101100111001101110111001001000111011101110000000001110111011001110000011101110100011101100110011101110111000001010001011101110111011101110111011100100111011101100111001100010001001101010111011100100101011101110111011101110010011100010111011101110100",
		"01110111011101110111001001110111011101110101001001100010011100100101010101110111011101110111011101110100011000000110000001100111000101110110010001110011011101110000011101110111011101110111011101100111011001000111011101110111011101110110011101010111011101110100010101110110010001100111011101110000000100110111000100000000001000010111010001110111011100110111011101100111001101110111011100100011011001110001011101110100011101010001011101110001001101110111011100010111011101110111011101110111011101110011010001110100",
		"01110111011100110111001101110111011101110111011101110010001000000001001100110010011101100111000101110101011100000111000001110111010001110111001001110011001000010111010101110101011000010111011100010111011101110111011101000000011101110111011101110111000101110010011101010111011101110000010100000111011101110111011100000011000101110101011101110110011101110001011101110111011101100001011101110111011101110001000001110110011100010011010101010001011101110111011101100101011101100011011101110110011001000111010001110010",
		"01110111011101110111000001110111001101110111011101110100011100000111011001110111011101110111011101110000001001110100011101000010011101010111011101110111010001110111010101110010011100100111011101110010010001000110011100110111010100100111011101100111010001110111011101010111011101110110011101110111011101110111011101110111000101000111011100100011011100110111011101110000011101110111001001110111011101010111010000000111001101100011011101000011011101110111011101110111000001110101011100110010011100000111010101110111",
		"01010001001101110010011101110111011101010111011100100111010101110111011101110000011100010111001101110010011001110111011100000100000000010111011101110111011101110111011101110111010101110111011101100111000101110111011100110111011101110111000001110101011000010100011100110101000101110111011101010000011100100110011101110111011101110111010101110111011101110111011100010111011100110111011101110111011101110111000001110010011101000000010001110111000001110111011101110111011101110100011100100110010100100110011101110000",
		"00010111011101110011011101110111001101000111011100000111000101110110000101110010000001110111000001100110011101110111001101110010011101110000010001110110000101110110011101010111011100000001001101110111011100100111011100110111010100100010011101110111011101110111011101110111010001110111001001110010011001110010011101110110011101100111010001010011011101110010000001110110011101110100010100010111010100010001011101110100010001110111011101110101011101110101011101110111000100010101011101100101000001110010011101110010",
		"01110000001101110111011100110111010001110101011100110111011101000111000101010111000001000111010101110001011101110111011101000111011100000111000101010111011101110111011100000001011101110111001001100011010100000111000100000011010101110101011101110111010001110110011100100010000101100001011101110111011101100111001001110100001101110111011101110101011101110111011100000000011100110111011100010111001101010100011101110111011101110111011101110100011101010011011101110110011101110101001000010110011101010111010101100001",
		"01110111011001000111000101110111011000010111010001110111011101110011001101110111001001000111010100100111011101110111011100000111010101110111011101110011010101110111011101110001010000010010001001110000011101110100011101110110011101010111010101000111001001110100001001110111011101110111011101110101000001110101011001110111001100100111011101010111011101110111011100000101011101010110001001000111011101110101011101110111011101110111000101000111001101010111011001010000011101110111011101110100011101100111001101100000",
		"00100100011100110111011100110000011101100111010001010011011001110111011101110111010000010111011101110111011100110111011101110111011101110110001101110111011101110111000101000111011101110010011101110001011101110001001000000111001101110111011101100011011100000111000101110110001101000111011101000111011101100111011100010111011101110111000000100111011101110111011100110111010100110110011101110011011101110100010001110001011100010111010100100111001000010010011100100010011101110111011101110111011101110110000101110001",
		"01110111011100010010011101000101011101110100010001110000011101110111011101110111011101110111011101110111011101110111011101110111011100000111001101110111001001110111000001110111011100010111011101110000011101110011011101110111011101110111011100110111011101110111010001110111011100000111001000000101011100110111010001110001011101110011011101100011011101000100011100100111001100100111001101010001011101010011011101110101000001110111010100110111001001110010000101110101011101000100010101110101001000100110011100100001",
		"01100111011101110001001001110001001100110111011101110111010000110111011101000101011101110110011101110111011100100110010001110111011101110111011101110111000101000001011101110111011101110101011101110111011101110001011101110010011101110111000100110111011101110111011101110100011101110001011101110111011100100111011000100111011101110101011001110001011000010111011101110111001001110011001101110111011101110111011101110111010001110111011101010111010101110111011101000000011101010111000101110111011101110010001001100111",
		"01110111011101110111000001110111001001000101010001110111001001110111011101010111011101110000001100110000001100110110011101110010011101110101011001000001000101110010011001110111011101110010011101110111001101000100011101110111011101110111011101110010011101010101011101110011011101100111011101110111000000000111011100110100000001010111011101110111011101110001011101110111011100110111011101110001011101110111001000110110010100110000011100000110011101110100011101110111001001000111001101110100011101110111011101110111",
		"01110000010000110101011001110111000101110100001001110111011100110011011101110101011101010111011101110111011101110111000001110111011101110111011101110111001101110111011100110010000000000111000101110011011100010111011101110111011101000110001101110011011101100010011101110111011001110111010101110111011101110001000100010111001000100111000001110111011101110110010001110001001000000011001001110111011101110010011101010111001001110100011101110111000100100111001101110100001001100111011101100111000101000111011101110000",
		"00010111011101110111011100010111000001110001011101100000011100010111010001110111011101110111000100000111001101110111011001110111010101110100001001110111010101110101000101110110010100100111010001110111011101110101001101110111000100010111010001110111011101000111001001110111011001110111001001110111001001110111011101110101000101110111010100110001011101110000010101110111011100100010011101110111001001110111011001110010011101110110011101000111000001110010011101110100011100110100011101110111010100100100011101110111",
		"00110011010101110001011101110111011101110001011101110111011101110111000101110010011101110001011101110111011101010000010101110111011101110111011100100111011101100001000001110111011101100111011101110111000101110011011101110111011101110111010001110111000100110111011101110010011101110101001101010111011101110001011101110111011101110111001101110111000001110111011101110111011101110111010000100111000101110100011101110011011100000100011101110011011101000111011101110111011101110111011101110111010001010000001100100101",
		"00010001011101110101011101110111011001010110011100000111011100100100000101110010000101110011011101110111001101010111001001110011011100010000011100010111011001110000011101000110011101000111001101010111011101110110011101110111001000100111011101110111000100100011000001000100011100010100001001110111011101110111001100100001011100110111011000110111000001110010001001110111011101100111011100010111011101110111011101110010011101100110001001010111011101110010011101110101011100010000011100110111011101010111001101110111",
		"01110111011101000110000100110111000101110111010001110111011100110011011101110110011101110111011100110100011001110111011101110010011100110111011101110001011101100111011101110101011101110111011101110111011100010111011101110010000101110000011101110111011101110000011101110111001001000110011101110001011001000001011101010000011101010111011101100111000101110011001101110010011101100111011101110110011101110101010100110100011101110111011001110111011101100000011001110111010000100111010001110111010101110111000001110111",
		"01110111011001010101011101110111011100100111011101110001011101110110011101100111011101100111011101110111000101110111011101110111011100100100011101110111011101110000011100010111011101110111011101100111011101110111011100010101011101110010011101110111011101110111010101110111011100100100011101110111011101110111010001110000011101110111000001110111010101110111001001110111001101110111001001110010011100010111011101000111001101000111010101110111011100100101000000100111001101110011011101000111011101110111000001110111",
		"01110111011101110110011101010011011101110101011101110111000101110111011101010111011101000010011101110111011100100011011101110110001101110111011101010111011101000111011101110010010100100111011101110111000101110111000101110111011101110010010100000111011101110111011100100111011100000111010101110001011101110111011101110110011101010111001001100111011101110101001001110110000100100111000101110111000100000111011101110111001001100101001001110111011101100110011100000111011100000111011001110111000001110000011100000111",
		"01110000011101110111011101110011011101100011001101110111000000010111000101010111000101110011011101110100011101110111010001110111000001110111011101110111010001110010011101110111011101110111001101110111011001110111011001110010011101110111001000010111011101100000010001000001011000100111011101100111011101110101010000000111001000000111010101110000011100000111011101110111001101000111001101110110011101110100001001110000010100100100000001110111000001110111011101010101011001110111000000010110000101100111011101110101",
		"01110101011101100110011101110111000000000111011101110110011101110111000001110111001001110111011101110111011101110111011100000000011101010111010000010111011101110111011101100100011101110000010101110111011001110011011101110111011100110111011101110101011101110001011101110010010101000011000101110111011101000111010001110111000000110100011101110111011101110111001000100111011100010001011100000010011101000101001100100111011100000111011101110111011001110001010100110111000001000111011101000111001000100010001101100111",
		"00000111011100010111011101110111011101110110010101100111011101100111011101110111011101110011011100000001011101110111011101110101011100100111011101010100011000010010011101110111011101110111011100110111011101110111011001000111001001110110011001000111010001110000001001110111011100000100011100000111011101110010011101110111010101110111010101110111011101100011011101110111011101110111001001110100011101110111001101110110011101000010011101110010011101110000011001000100001101110100011101110110001000100111011100010010",
		"00100111010001010111011100010010000000100011011101100111011101100111010100100111011101000001011101110000010101010111011101010111000101010111011101110111001101110000011101110111001101110111000101110110011101010011011101110111011101110101001001000001000100110111011100010011011101100111011101110100011100000111011100110011001101110111011001110111011101110100011100010111011000010010011101100111011100100111010101110111011101000111011101110111011100100010000100010111011001110111011101110010011101110111011101110111",
		"00100111011101110111011101110111000101110111011101010111011101000111011100000000011101110111000100110110001001010110010001110001011100010111001001110111010000110100011101110010011101110010011100110111011100010010010101110111000100000011011101110111011101110111001100010000011101110111011100000111001100000111011100000101011101110111010001110111000101110111011101110111010101110000011101110111011101110111011100110001000101110111011101110111011101000111000001100001011100010111011101110000000001110111011100100100",
		"00110111011000010111011001000111010100100101011100000111000101110111011101110101001001110100011101110111011101110001011101110001011101110111011101110111011101110100011101110110010001110111001101110010000101010111011101110111010000100111011001110111011101000111011001110111011100100111000001110111011100010101011101110111010100010111001101110011011101110111011101010101011101110111011101110011011100010010001101110111000101110111011101000111011101010111011101110111010000000111010101100111011101110010011101110011",
		"00010111010101110010011100100010001101110110001001110011001001110001000001110111011100100101010000100010011101110111011100110111011100010000011101110111001101000000011101110111011101110101000101110110011100110010010101110111011100000011001101110111011101110111011100110001011101110101001000100111010000010111010101110011011101000000011100100100011001110111011100100111011101110100010101110000011001000111010101000111011001110111011101110111011101110111000001110111000001000111011100000111011101110111001100100111",
		"01110011011101000010011101010110000100110111011100000111011101110110011101110111011101110001010001110111011101110111011101110111011101110111011101110111010101110111000101000111000101110100000001110101011100110111001001100011011101010111010000010111010100100100011100000111011100110111011101110111011101110100011101110111010101100111001100100111011101010010010001110101010100010111011100000111000100110010001001110111011101000100011101110011001001100111000000010111000101110111011101100111011001110111000101110111",
		"00110111011101110000011100010111001000000111011100010111011101100111000100110001011101110111011101000111011100010111011101110110011101100111011101110010001101110111010100100111011100010111011000110111011100010110011100110111001001110001011100100111000001110111001001110111000101110111001100110111011101110111011101000111011101010111011100010111010101110100011101110111001100010111011101110001011100010010011101110111010000000111010000100011011101000101011101110111011101110001011101110111011001110011001101110111",
		"01110110011101110110000001010111011101110111011101110011011001110111010101110111011101100111010101110100011001110111011101100101001101110100011101010011011001110111000001110111011101110111011101010111011101110001011101110101011000100100011101010111001101110111011101110111011101110111000001100111000100110100011100110110011101110111011100000111011101110111011101110110000100010111000001110111000000010001011101110101010001110111011101110111011100010111011101100111011101010011000101000111011101110100011100100111",
		"00010111011101110001011101110111011101110111011101110100011001110100011101000000011101110000010001110110011101110111000001110111010001110011011101110111000000100101011101100111001101110111001100000111010101010111011100010111001101110010011100100111010101110111011101100111011101110011011101110110001000100111011100110111001000100111000001110111011100100111011101100000011100110111010001100100010001110100011100010111011000100010011101110111010001000001011100110001000100010111011101110100011101110110001101110111",
		"01100000011101110011011101000111011101110000011101110111011101110111011001110000011001110111001101110011010001110111011100110111001001100111011101110111011100000111011100010111011101110111000001000000001001110011001101110111011101110011011101110101011101010111011101110111000001110111011101110111011101110111001100010111001101100111010100100101011101110111011101110111011100010111011101110111011101110111011101110111011101110100011101000100000001010011011101110111001101110111011101110111011101110101011101110111",
		"01110101010101000111010000000110000101110111010101110011011100010010011101110010001101110111001101110001001101110100000101100111011101110100001100110111011101010111010100110000011101110000011101110111011100010000001101000110000100000001011101110101011000010111001001110111010001110110000101000000000101110111011101010100011101110111001001010111011101110000001101110110010101110101011000100100011100000111011101110101011101000111011100100010011100000000011101110111011101110111011100010111010001110111011100000111",
		"01110111011101110111000001110111000001110111011100010111011101010010001101110001011101110111011100010111011100000111011001110101011101110111011001110010011101100111011000100000011100010111011101110110000001110111011101110111011101110111000000100010011101110111011101010101000001010111010001110111011101110111011001110000011101110111010100010111011101110111010001010100011001110111011101110111001100010111011100110001001101010001000100000110000101110110011100000001011101110111011101110111010000010010000001000111",
		"01110111011101100111011101110011000100000111000001110111011101110111011101110111011101110011011101110111011001110111010100000100011100110111000101100111001101110111011100010111010101110010011101110101011101100110011000010111001001110000011101110010011100010111011101110111011101110011000001010111011101000000011101110111001001110101011101010111001001100111011001110110000000010000011101110111011101110000011001110100011100110111011101110111011101110111001000100100010001010111011100010111011001110111011101110110",
		"01110101011100010001001101110010011100110110010001110111011100100111000101110111011001110111010101110111011101110111011101110111011101010110011101010110010101110001011100110100010100000011010101110100011101110111011101110111011001110010011101110010011000110111011001110000011001110111000001100001011100100111000001110001011101110111011100100111011100100111011100100111001001110111011101000111011101110111010101100111010001110111011101110111010101110110011101110111011101110111010001110100000101100001001101000001",
		"01010010011101010111001100000000011101110111011101110100011101110111001100110111011101110111010101000111011101000111011001110111001101100111011101110111010000000111010001110111010001110111001101010110011101000111011101110111011101110000011100000111011100010100011101110000011101110011011101110111011101110000010000000011011101110001000001110100011001110111011101110110011100100110011100000000011101100111000001110111011101110111011100010111011001110110000101110011011101110101011101110111011100110110011101110111",
		"01110111010001110111000100010111011101110111001001110101011100010010010101110111011000010111011101110111000001100111011101110111000101000111001001100101011101110000011100110111010000000111011101110111000001110001010101110111011100010111011101110111011101110111011101110111001101110100011101110000000001100111010001000001011101110111011101110111010000100101010000100010011001100000011101110111011101110001011101110111011100000000011101110010000001110111011100110111001001110101011101110111011101000111011101010111",
		"01000111011100110111010001000011000101110111011101010111010001110101000101110111011101110111000101110101011100100100011101110111001101110010011101110011000000010111011101000111011100010111011101110111010001100010011001110101000000000111011101110111010100110111011101000011000100010111011101110111011100100111001001100111011100100110011101100111011101110001011101110111010101110100000000100110011101110111000101110111011101110011011101110111001101110111011101110111011100010011011101110111011101010000010000010111",
		"00010011010101110111011001110111000001110111011001110010011100110101000001110111011100100101011101110111010001110111011001110101001101010110000001110101011101110111011101110111001100110111010001110111011101110111011001110001011100000000011101110111011100000111011101110111011101110010011100000101011100100001010001110111011101110111011100000111011101000010011101110010010101110111001101100001010100010111011101110111010001110111001001110001011000110111001101110111011100010111011101110111011101110100011101110111",
		"01110011010001110111000001110111000101110111011100100111011101110111000000010110011101010111010100110111011100100111000100110111000101110011010001110111011101110111000100010000011101110111011100100111011101110010011101000100011100100111010100010000000101110000011101110000011101010000011001000111011100100111010001110100011101110010000101110111011101010000001101110111010101110111011101000111000101100000010000100010011101000111000101110111011101110110011101110010000001110111010001010111010001110111001001100111",
		"01110100011100000111001001110100011101110010000001000110011101110000011100100111010101110110011101110111001100100111000001110010010101110111011101000111011101000010011101110111011100100000000000100100011101110111011100100100011001100010000100000110000001110011001101100111000101110111011101110100000101110111010101110111010100010110011101110001011101110001000001110111010001100111000001110111011101000111011100110111011101110010011101110111011101000011011101110100000001110101000101110111011101110100011001000111",
		"00000010011100010100011101100001011101110011010100110100000100000111011100100111011101110111011101110010011100010111010001110100011101000111011101110111011101110111011101110111011100110000001101110101000001000111011100100111000001110011011101000111001101110111011100110111011100100111011101110001011100100111011100100111011101110010011101110000011101110111011101110101011101110111011001110001011101110011011100010111000001110100011001110111011001110111000001110111011101110010011101110111011100100111000001110011",
		"01110111011101110101010101010111011100110101001100000010011101110111000101110111011100100111001001110001000000100011011101110111010100000011000101110111001001010111000101010001011100010101011101110111011100100111000001110000010000100100000001010111001101110111011101010011011001000111011101110111011101100111011100100111011101110100011101110001011100100111011101010111011100000111011101110111011101100101011101110111011101010111011000010111010001110111011100000111001100010111011001110100010100110100011100110111",
		"01110011011100010111001001110011001101110111011100010111000101110010011100100011000000100111011101110011011101110111010101000110011101110100000101110111011100010101011101110001011100010111010001110111011101110010011101110111011101110100011101100111001101000010000101110111011001110111011100100111000101100100000001110111011100100011011101110111011001110000001101110111001001110111011101010011011101110100011101100111011101110111011101110101011100000111011001110111000001110111011100100111011100110001011100100111",
		"01000000011100100001011101100001010000110111011101110001010100000100011101110001011101110000011101100000010101110111011101110000011101110101011100010111011101110111011100100111011100010111011101110111011101110111011101110111000101110001011001110111011101010111001001110000011101110111011001110010011100010110000101110111011101010010011100100111000000110111010000110111011001110010010101110111001000100001001100100111011101010011011100100001000100000101001101110011011101000111011100100011011100000111011101110000",
		"00010000011101110101011100000111011101010111011100010111011100110111001001110111011100110101011101110111010101110100010101010111001001110111011100110111011101010111010100010111011100110100010001110110001101110111010001110111011101010111011101110001010100000001011101010111011101100001000001000001011101110111011100110110001101110111000100110111011101110111010001110111011101110111011101110111011001110111011001000101011101110011011101110111011001110111011101010111001101110010011101110111011101110111010001110111",
		"01110111011101010111011100110010011101110111011101110110011101110111011101110110000000000111011101100101001001110000011101010011011100110000000001110111011100100001000101010111011101110000011101110111011000010100011101110111011100100111001000010101011101110111010101110100001101110111010100010111011100000101000100110110011101110111011000100111010101110100010001110111011001110011011101110111011100110011000000100111000001110101011101110111011101110011011101110111001001100101011101110111001100110111010001000111",
		"01110111001100100101011101110010011100110010000101010101011101110010000100110111011101110111011100100001011100110000001101110101011101110001011101110011011101110111001001110000001101110100011001110111011101010101011101110110011100100111011101110101011101110010011101110111001000000101011101110110011100010011011101110111011100000111011101110111011101110100011101110010011001110000011101110111011000010010000101110111011101110110011101010111011100010110011101110011001001110111011101110010011101110111011101110101",
		"01110111000100010111011101110111001101100100001101000111001001110111011100110001011101110101011101110111011101110111011101010111010000110111011001110111011100110101011100110111011101110111010101100111001001110100010000000111010001110010011101110111000001110010001101110111010001010111011101100001011101110100011100000111011101110001011101110111010101110111011101000111001101110111010001110011010100100111011101110111011101110011001000100111011101110111011100010111010101100010011100000100011001110111011100100010",
		"01110100011100000110010101110111001001000111011100010111011101110101011101110010011101110111011101100111001101110111011101000010011101100111011001110101001101100111011101110010011101110111010001110111000101110110001001110111011101100001011100000000010001110111011101010111000001110111011100010111011100010100011000100010000100000111011101110011011101110001011000000110001001110101011001110111011101110101011101000011000101110111010100110111011100000111011101110001011100110110001001110111001101110111011100010111",
		"01010111011101110111011101110111000101110111001001100111001001110010000101110111000000010010011101110100001001110111011001110111010101110111001101110100011101110010000101110010011100000111011100100111000001000111011101110101010101110111011100110111011101100111011101000111011101010111000001000100011101110001011100110000000001010000011101110111011101110000011101110111000101010111011101110111000101110011011101110001011100100111011101000111001001110110011101100111010100110001011101110111011101110111001100100011",
		"01110101011101110000011101110111011100000011010100010010001001010100011001000101011100000011011101100001011100100100011101000100001101110111011101110111011101100111011101000110011000110101011101110111011101110110011101110100001001110001010100100101011101110000001000000111011101110111011101110111010000110100010001100010000101110111010001110111011101110111011101000111011101110001010101110111010001110111011101110101011101010111001100110100011000010110011101110000011101110111011101000111011101010000000101110111",
		"01110111010101110111011101110000001001110101010001110111010100110111011101000111011100100101000001110111011101110010011101110001010001110010011101000111011001000111011101110111001000000011011101110111011101110111000101110100011101110110011101110000000101110000010101100001000101010000011101110111011101110111011100110111000101110100000001110000011101110111011100110100011101110111010001110111011100010111011101110111011101110111011101110111011101110111010001000111011100010111011100100011010101110111011101110111",
		"01110111011101010111011100010111010101110111011100110111001000100001011101110111011101110101011101110000000001110101011001110101000101100111011101000111000101110000011100100011000000010000011101110001011101110111011100110111001000100110011101010111011100010110010001110111011101100010011100110001011000010100011101110000011100010111011101110111011101010011011101110111011100100110011101110111011000100101011101110111011101110011000000100010000101010111011100000001011101110100000001010111000001110111000001110111",
		"01110111000100010010000001000111010001110010011000100111011101110111011000110111011101110111011101100001001000110111011001110000001001010010001101110111011001110111010101110000011101110110011101110111011100100010011100000111011101110111011101110111011101110111001001110101011101000010010000110010010001110110001001100111011101110111011101010100010101110101000000110101011100000010010001110000011100000000011101110001001000010111000101110111000001110111001000010110010101010111001001110011010001110111011101100111",
		"01110111011100100111011001110111000000100011010101100011001101110101011101110100011101000101011101110111000000010111011101110111011101110111001101110111011101110111011101110111010001110100011001110101011101110000011100110001011101000100011100100100010101110110001001000111011100000101000101110011011101110111011101110111011101110111011100000111011101000111011100110111011001110111011000110011000101110110010101110110001100100111011001110111011101110111010001110010011101110111011000110111011101110111011101110000",
		"00010111001001110011011101110111011100010111011101110111011101110100011100100010001101110010011101010100011101110011011101110111011101110111011101000011011100010111001101100111001100100101000000000011011001110001011000010011011001110011011101000111011101110101011101110111010101110111011101110100011101110010000000110001011101010111011101110111011100110111011101110001011101110111000001100101011101110001011101110111011101110111011101110111001000100111011101110111011101000110001000110011000101100101011101110101",
		"01110111010101000111011101110001011100100111011101000100000001100111000101110001001000110100001000000111011101000100011101110001011101110111010001110100010001110111011101110101000000110111000001110011011101110111000001010101000101100000011101100101011101110111011000110010001001110000011000100111000100000111011101110101001001100111000101110100011101110110001101110111000100010000011101110011011101100010011101110111011101110111000100010101011101110101010101110011010001110100011101110111011101010111011101110110",
		"01110001011100010000011101010111010001110111011101110011011101110100000101110111011101110000001000100111011101110111001001110110000001110000001000110011000001110111000001110111011101110101011101110011010000010111001100010001011101100111011101100001011001110011011101110111011001110111011101110111011101110111001101100111001001110000011101110111000101110111010001110111011100000111011101010111011101110111000001110011000100100111011100110111011101110111000000100111001001110111011101100010011101110111011101110111",
		"01110111010100110111011101010010011101110111011100110110011101110111011100100000011001110111011101110111011101110111011001010111011101110111010001110111000001010111010100110111011100000111011101110001011001100100001001100111010101110111011100000010011100010111011001110111011101100001010001110011001101110101011101110111010001110000011101110111011101110000011101010111011100000111000100100000011100010011010101010110011101110101011101000111011101110111011001110111001000010111011101110111001101110010011100010110",
		"00010010011001110111011101110111010101100111011101110000001100010011011101110111011101110101011101000110011101110111011101110111011101110111011101010110001000100110000000110111001101110111011001100111010101110111011101110000011100100100011100110111011100010000000001110111011000000110011101110101011101100100000000110011011101000101010101010100010101110111011000010000001001110001011001110111000001110111011101110111001101110111011101110011011101110010011101110000011100000111011101010111001101110111010101110100",
		"01110111011101110111010101100110011101000000011101000110000101100000001001110001011100100011011100100000011100100111011101110111000001110111011001110001010101110111001001110100010101110001001100000111000000000000011101110010001001110001011101100111011101110111000001110111011101100111000101010111000000110011011100110111011101010111000000110111011101110111001000000111011101110111011101110111011100110111001001110100011101100111011001110101011001000111001001110101000101110111000100100100011001110111011100000001",
		"01000110011101100010000101110111011101110111011101110010011101110111010101110010011100010101011101110011011101110111011101110000011101110000011101110110011100100111011101110010001001110111011101110110011001000111010100010001010000110111011101110011011101110111011101110001011100110111000001110000011101110111010000010001001101110001011100010010001101110111011101100111001101110111011101110111011100010111001101110111011100010111011101010111010100110111010101000011011101110000011101000111011100100100010001110111",
		"00010111011000010111011101110111011101110111000100000111011101000111001100100111011100010111010001000111000101110010010101110000010101110110011101110000000101110010011100000000001001010101011101010111011101010111000000010111011101110010000001100011001001110111011101110111011001110001010100010011010001110101001001110111011101110011011101110101011101110111010001110110000001110111011101110111011101100111011101110111001001110100011101110111011100100111011101110111010101000011011100000101011100100110010101110011",
		"01110001011101110111011101110111011101110011000001110010011100110111011001000111011101010111011101110111011101000010011100100111011001100111001101110101010101110111011100100111010001110111011100110111011101110111011101110111011001110111011100000111010001110000001001110111011101000111000100110111010100000111000000110111011101010110011101110111011100010111011101110111011101100111011101010111011001100111011101100111001101110001000001110111001001110011011101100010010101110111011101010011011100000111011100100111",
		"01110011001101110111001101110111011101000111011101110000011101000111011101100111011101110111010101110111000101110111001001110111011101000111000000010111011101110110010001110101010101110111001001010100001001110000010100010111011101010101011101110111011101110100011101110111010001110111011100110111011101110100000101110000000000110001001001110110001001110000000100110111000101010001011100110100001100010111000101100111011101010000010101110111001001110010011100000111011100100111000101110111010101100000011101110100",
		"01000111010101110100011101110111001001110001000101110111010000100101001101110111011101110111001000100010011101110100011100110001010101110100011101010010011101110100010101110111011101110111011101110111001000000100010101010001011100000111000101110111011101110010011001000100011101110000000101000111010001110111011100100111001101110111010101100100001001110010010101110111011101100010011100000100011101110010010100110111011101110111011100010111010101010111011101100111011101110111011101110011011101110100010101110110",
		"01110111011101110101000101110111011101100111011101010111001001110111011101110111011101110000011101110010011101110011011001110111010101010111011101110111011101110111001001110010011100100000011100000111010101110111010001110111010101110111011101010100011001110111000101110111011100000111011101000100010101110001000001110100001101110111011101110010011101110111011101110111011100000101001001000101010001000111011101110001010000010110010101110111010001110111011101100010011101110110011100110110000000100010011100010001",
		"01110111011100100111000101110101001001110010000001000111011101100111011100010100011101110010011101110001010000100111011101110111011101110111011101110011011101110010011101110111011101110110011100100111011101110111011101110111001101110000010001110010011100000111011101110101000001110111000000000001011101010101000001100111010001110001011101110111010001110100011101110111000001100111011100100111011101110101011101110111011101110111011101100111011100010111011100100001000101110100011100010111011100110110011101010111",
		"01000011011101000111001001000111010001110000011100100111011101110111000001110010011001110011011100100111010100110111010000110111011101100101011101110010011101110111010101110111011100110001011001010100011101110011011100100101011000000001011100110111000001110111011101110111011101110111000001110110011001100111011100110111010100010111011101110101001100000100011101110111011100000111001001000111000001110111011101110111001001110111011100010110010001110111011100010111011100100111011101110100001101110011011100010111",
		"01110100000101000101011101100111011100010101011101110111001001110111000101110010011100100111011101110101001001110011011101110111011101110111011101110101010100000111010101000111010101010111011101110001010101110111011101110111011101110111011101110111011101110111010001110001011101110111011101100111011101110111011001010010011101000111010100100111011100000111011100000101001101110001011101110111000101110101011101000111011101100111011100010111011101110110011101010111011001110101001000100111010001110111011001110111",
		"01110110000101110000011101110111011101110101010001110111010101010000011101110111011101000111011101010100001101110101011101110110011101110111011001110111011100100110011101110001011100100010001100100111010101110111001001110000011101110001011100010111010001110111011100000111010101110111011000010111011101110111011101110110001001110111010000000001011101110100011101110111000100110111011101110111011101110111011101110111011101110001010001110111000001110111011100100111011101110111010101110000000101010010000100000111",
		"00010111011101110101011101100111011101110111011101110010011001110001011101100111011101110111011101010111011101110111000101110111011100100111010001100010010001100111001101110001011100000010011101110111010001110001011101110111011101110110011001110001000101110111011101110111011101010010011101110000001001100110011101010111011100100111010100010111001001110111011100000111011100000111011101010111011101110111000001110011011101010111011100010011011101110010011100100100010100100111001000110111011101110111001000000111",
		"01110101011101110111010101110110010000100111001001110111011101110000011101110111011101110111010001010111011100010100001001110011011101110101011101110111011101110000000001110111011101110110011101110111010101110110011101110101000000010111000001110011011101110111011101110010001001110111011101110111011101110111000101110111010100000111001001110110011000000011010101110000000101110111001101110111011101110111000001110111011100100111010001000010011101000111010100110111001101110111011101110110000000000111000000000111",
		"00000100011101110111001001110111000100000111011101110011010001110111011100010111010101010111010001110111011101110011011101110111011101110111011101110100011101110100001001110101010100110000011101110011001100110111011101110110011100100100010101110011001001010111011101110111011101110111011100100111011100000001011101110100011101110010011101110111001100010111011101110111001001110111011100000111010001110111011101110111011101100111000001110111010100100111011101010111011100100111010001000111000101110111001001110101",
		"01010111011100100101011100000111011001110111011101010010010001110010010001110111011101110101001000000111011101110010001101110000011100110111011101110111011101000111011001110000010001000101011101110001001101010111011100000111011101110110010000010100011101110111011101000111011101010111011001010111011101110111011100010111011100010010010000010111001101110111011101110111000101110111011100100111011101100111011000100100011001110111001001100001010100010111010000110111011100110110011001110010011001010111011101110111",
		"00000111011101110010001101110111010101110111011101100011011101100111011100110011010101110111011101110111001101110100011100100111000101110111000001000111011100100111001101110000011100010111000001110111000000110000011000000000011101100111001001010111011100010010011100110111011100000101011100000111011101110110011100110111011101110111000101110000011101110111001001110111000101110111010101110111001001110100011100010110011100010010001001110111011101110111011100110101011001110111011101110001011101100111011101110111",
		"01110110011101110111000101110100000001110111000001110000001101110101011100110111011001110111000000000011011101000111011101000111011101110100011100000010011101110111010101110111001101110011011101110111011101010111011101000011001000100100011101000111011100100110000101110111001101110111000101000000000101000110000001110100011101010001000101110111011101110011011101110001011101110111011101000000001001010000011101110110010001110111011100010100011101110111010101110011011101110111000101110010010000000101000001110011",
		"01110111011001110101000101110111011101110111001100010111011001110000011001110011011101110111011101000111011100010101000101000111011100110111000000100111010001110011010100110111000100100111001001110111011001110111001101110111011101110111011101110111011101110011001001110001011101110100011101110111011101110110011101010010010100000110011100100100011101110010011100100011010101110111011101100110011100010011011100100010010101110111010101000100010001110111000001110111001100010010011101000111010101110111011101100100",
		"00110001001001110111011101110111011101110111001100100110000101010111011000100111011001110011000001110111001001110111000100000111011000110111011101110100011101100111011100010111011101100000000100010111000101110001010100100111011101010111011100000110011101100011011100010111011101110110001001110111011100110111000100110110010000110011000001110000000101100111011101110111000000110101011100110111011101110101011100000111011101110000011100010011011001110111001101110111001101110111011100110111011101110000000001000111",
		"00100111011001010111011001100111001001100111001101110111011101110111011101010111011100010111011101110111011101110111011100110111011100010111001001110001011101110111000001110000010100100111011101110111011101110111011101110111011100110110000000100111010001010111010101100010001100110000011100100111011100010100011101010111011001000101001101110111001101000110010101100111000001100111011101110011011001110010000001110010010101010110011101110111011101110111011101110111011101110011001001110101011101110111001001110000",
		"01110111011100000111011101000111011001110111011100110110011101110111011100010111011101100010011001100111000101110111010000110111000001110111000001110111011101110110011100000010011101110111011100100111011001110110011101110111001001110010001100110111011101010101011100100111011101010111011101110100011100100100001000110100011101110100001001110111011101110011011101110001011100010111000100100001011101110111011101110111000100110111011101110111011100000000011101110111010100010110010001110111011001000111011001110110",
		"01110111011101110100000100100001011100110001011001000010011100100111011101000111010101110011011101000001011101000100011001110111011101110110010001110111011101010001011101110111011101110111010001110110001001010110011101110000001101110100011101110111011101010111011101110110011101110111011101000001000001110110010100100011000101110111010100100111001001000111000100110100000000100010011100000111001101110101011100000111000001010000010000110011011101110110001101110111011101100111011101110001011100010000011101110110",
		"00110111001100010100011100110111001000100111011001110111010101110011011100010001011100110011010001110111011100010111010100100110011101100111010001110111011101110100000101110111001001110111011100000011011100010011001001110111001101110010000001000100010101110111010001110111011001000111000100100111011101110110011101110011010101110111011100100111011101110011011101110111010001110000001000100100010100100111010001110010011101110111011101100111011101110111011000010011001100010111011101010000010000010111011100000111",
		"01010111011101110101011101000011011001110111011101010111011001110111011100010010011101010001010100110111000001100111011101000111010001110111000000110110011101110111011101000101011101110111011100000111011101110101011101110111011101100111001100100110011101110111011100000111011101110111001001110111011100100111000000100100011101110000011001110100011101000111011000110111001101110111011001100101010100100111011101110111000001100111010100010111011101000101001001010111011100000000011000100111001000110011010101110111",
		"01000010011100000111000000010111000100100101010101110111011101110111011100000100011101110111001001010011001001110111011101110111011101110010011101110111010001110001011101100111011100110101010101110000011100100111011101110110011101110100011100000111010000000011010001110111001000000101011100100111011101110111011101000011001001110111011100100001001001110111011101110001000001110101011101110101011101110111011100000111000101010111010000010011011101110110011101110111011101100111001100000111001101110111000100110111",
		"01110111011101110101000001110111011101100111011101100111010001110100011001100111011101110100000001100001011100110101000101110010001101110111001101110111000001110011011001000110000000110101000001110111010101110111011101110110011101110100011101110110001001110111011100000001011101110111011101100111011100010000011000000111010101110111001100100111001001110111011101110111011101110111010101110111010100000111001001110111000101110101011100110111011100010111011101110010011101110101011101110101000101110100001001110111",
		"01110001010001110110010000000101011100110010011101110100011101110111011100000111000000010111011101110111011101110111010101110111011101000111011101110010011001010111011101100111011101110010011101110010011101110111010000110110000100000100000100010111011101110111000101110110010100110111010100010111011101110111011101110110010001100111011101110010000101110111000101110100000100100111011101100101011101110111001101110111001101110010011101110001010000110111011001110111001001100111011101110101011100010111011101010101",
		"01110011011101110111011101110111011101110111011101110111011101110011011101110111011101110011011100110111011101110111011101110111011101100010011101110011000101000011011101110111001001110111011101110101011101110111010001110010001000010111011101110101011101110001011101110111011101100111010101100100011101110111000101110111000001110100011001110111010000110111011100110111011101110111011101100111001101000001011101110000011101100111011101010011001101110001010001110111011101110101011101110001001100000100001101110000",
		"01110101011101110111010000110111011101110111011101110111010100000100001000000111011000100111001001110111011101110111011100110111001100000111011101100111010101010001011101110111011101100011011100110101011100110000011101110111001100000111011101110111000000000111000001000111011101110111010101110111011001110111011101110111011100000011011001110100010001110010000101110011011100000111011100100111001001110111010101110111011101110111011001110101000101110111010100000111001001110111011100100111010001110111011101100011",
		"01110111011101110111011101110101010101110100011001110001001100110111011100010110011101110111011001100111011001110111010001010110011101110111010000110100011100100111010100000110011101110110000100100111011100100111010001110000011101010111000101110111011101110111011101110111011101110111011101110111011101110111011101110011001000100111011101110111011101110000000101110111011100000111001101110111011101110111011100000100011101110000001101110010011101110111000001110111001101110011011101110010000000000001011101110101",
		"01110010001001110110011001110101011101110001000001110011000000100111000101110111000000100111011101110101011001110010011101110111000000000000011001110011011101100100000101110110000001110111001101110111000100010111011101110111011101100111011101110101011101110100000100000111010001110110011100100111011100100111001101110111011101010000001001110110011101110101011101100111010101110111011101110110011000010111010001110111011100000111011101110100011100010111001001110110001000010111010101110000011100100010011100100111",
		"00110111001100000111011101110011010001110111001000110001011101110111011101110011011101110111011001110001011101010111000100100101010001100111010100010111000000000111011101110111000001110111011101110110011101110111011100100111011101110111011101100111001001110110011100000111011101110011011101110111001001110111011101000101011101110000001100110111011101100111011101010111011001110111011101110000000001110111001000110011011101000111001001000111011100010111000101110111011101110111000101110111011101110111000101110010",
		"00000111011101110111011101000111000101110111011101110111011101000001011100110111010101110100011101110111011101100111011100000111011100010111011101110011011101110111001001110111000001110111010001110111011100100100011001010111010001110101010101110000000100000111010101110101011100010010010001110111000101110111011101110111001001010111011100100011000101110111010101100101001001110010011101110111011100100001011100010111011101110111011100010111011101110001011001110111000101110111011100010000011101000111011101000011",
		"01110110011100100110011100000101001100110001011101110011011101110001011001110101011101110111011101110000011101110111011100010010011101110110011101010111001100100011011101110111011101100111011101110111000001110100010100110111011101110011011101110111000100000111011101010001000001110001011100100111011101000111011101110111011101110111011100000111011101110111011101010111011100010111011101110111011101110111011101100111011101000011011101110001000101110111000101110111001001110111011101110111000001110111010101100111",
		"00110111011100110000000001110111001100100100011101110111010100000111000100100111011101110101011101100111001000100111011100000111011101110101011101110111010100110101011101110111000001110111011101110010011100100100001100010111011101000101011101100011011101100111000101110011011101110010011101110000000101110010011101110111010001110111011101110000011101110111000000110111011100000111010101000001011101010111000001110100000101110010011100110111001001110111001100000110011101110110011100010111011101110111011101000111",
		"00000001011101110110010100100000001000000101011101110111011101110101001001110111010000010010011101000111001101110111011001010011011101110000001101110110011101110100000101110111010001110111010101110101010001110111011101110111011101110110011101110111011101110111011101110111011001110111011100100111001001110000011001010000011101100010011101110111001101110111011101110111010101110111011100000111011101010101011101000011000000100111001101110011011001110001010000110111011101110111000001110111010001000111001001110011",
		"01110111011101110111001001110111011100010111011101110110011101110000011101100111011101110111010001110111011101110011011101110111011100110111010101110111010000100111011100000011011001110111011101110111011101110001011101110111011101110010011101110100010101110111011101110111011101110101001101110101011101110010000101100010011101010001011100100001011001110111011000110011010101110111001101110111001000110101001100000111011100000111010101110010000100010101011101110110011101110111011101110111011100100001001001110001",
		"01110111011001110101011101100111011101110010011101110111011101110111011101110111011101110111011101110111011101110010011101110111011101000111001001110110001001000111011101110111011101110010011101110111011100100111011101110000010001110111001000010001000101110111011000010110010000000010001001110010010101110010010101110111011101110111011101110010001001110000000000010011011101100111011001110101011101110111011101000100011001110101000101010011011100100111011100000111011000100001011101010111011100010001011100000111",
		"01110001010101110000001001110111011101110111010001000111000001110111000100110100000001110111011000000101011101110111001101110111011101010010001001110111011101110111011101100111011101110111011101110000011001010111010001110111010101000110011000000000011101110101011100100101011101110111011101110011000101110111011101110001010101000011001001110101011001110001011100000111011100110100011101000010000101110111011101110111011100010010011101100111000001110011011001110000011101110001001001110110010001110111010101110010",
		"00100010011101110111011001000111011101110111011100010111011101110101000001110111011101000111001001110111011101110111001100110011000101110111011100100110011101110111001000000111011101110111011001010111011001100111011101010111001101110110011101110101000100100111011101110111011101110111011000010111011101110111000001110010000000000111011101010111011100010111010001110111011100100111011101110111011101110111011101110111001101110011011100110111011001110101011101110111010000100000010100110111011101010110011101110111",
		"01110010011101110101011101100111011101110111011100010111010100010111010101110111010000010101011101110111011101110101011100100111000001100111011101110111011100010111011101110111011101110111011101010111001100000111010101110111010001100111011101110101000000100111011101110111011101010101001100100001011101000111011001000000011100100110010000110111001000000111001001110111000000110111011101110111011101110111001101010101000101110111001101110101010101110010010001110100011100000000001101110111011101110111011001110001",
		"01000010011101110111001100010000011101110101010101110000011101010100011100110110011101110101001001110000011001110000011100000111011100000111011101110111010101100111011101110111010001110111011100100110000101110111011100010010011101110111000100110110010001110111011101110011011101110111011100100111011101110101011101110101010100000111000101000111011101110111010101110111001101110101011100110111011101110111011101110111011101110001011101000000011101110110001000100100011101110111011000000111011100000111011101110111",
		"01100111010101000111010001110101011101110111011100000001011101110111011100000110011101110111001100110100011101110111001101110101011100010111011101110111011101110100011101110011011101110011010001110111010100000001010000000111011001100011010001110111011101110111011101110111011101110111011101110100011000100110011101110011011000100111000001110111001100000111011101110111000001110111011101100110011101110000011101110111001000000111001100010100011101110111010100000111001001110111011101110111011101110111011101110111",
		"00110111000001110110011100010110000101110111011101110111011101110111011101110111011101110100011001110100011101110101001001110111000100110011001001010111011101110111011101110111011101110100011101110011001101110110010101110111011100100111001000110101011100000111000001110010011100010111011101110001011101110111011100010010001000010111010101110111011101110111011101110111011101000111011100010000011101110111011101010111011101110100001001110111001001110111000001110100000100000111011101110111011100010111001001110001",
		"00100011011101110011011101110101000001110000011001000111001001110111010101110111011100110111000001110001011101110100001101110111010101110111001001010111011101110111010001110111010001110000000101110000011101110111010000100111000100000000001101110111010001110011011101110111011101110111011101110110011100110111011100100111011101110111011101110011010000000000011101100111011101110001000101110111011100100111010001110101001100010111011101110111001101110111011101110010011101110001001100100101010001110111011101110111",
		"01110111011000010111011101110011011101110111000000110000001100100000011101110111011101110101011101110111001000010111010101110101011101010111000100100111011100010011011101110111011101110110011101110111011101110101011100010111011101010010011101110111000001110111001001110111011101110001010000010111011100100011011100110111011101110111011101110101010000000111001000110111000001110111011100110111011101110000011101100110011101100111011101110111011101100111011000110101001001110001011101100111011101110111011101110001",
		"00110111011101110000010001110111011101110100010001110111010001110010011101110111011101110011010100100011001001110111011100010111011100000001011101100100011101110111001001110100011100100110001000010011011101110111011101110000011101110110001001100010011001110111011101110111011101110011010000010101011001110011011100000111011001100100010001110111000101110111011101100111001001110111000101110111011101110000011101110111010001110000011101110000011100110111000101110000011100000001011101100111000001110111001001010111",
		"00110000011101000111011101110110011101000111001100000000001100110101010000000111011001010111001001000111010101110111011101110111011100000111011101110111011101110100010101110000011101110100011101110101011101110111011100000111011001110111011101110111000100100111011001110001011101110111011000100111011101000101011101110111011100010000011000100111000101010111001100010000001001110111011101110111001101110111001000100111001100100111001101110111001001110101001100010111011101110010010101110001001001110110011101110000",
		"01110111010000110111011100000111011100100111000100000000011100010111011101110100011001110111011001110111011001110111011100100111011101110111000000010111001101100010011100010100010100100111010001110011011101000010001100110111011101110111011101110000011001110111010101110001010100110011001101100111011100000111010100100111001001110100011100000111011100100111011101110111011101110001001000010101000000010010000001110011001101110000000101110111011001110101011101100111010101110111010100010011010001110111001101110111",
		"01010001011101100000011101110111010001110001000100110111011001110111001101110011001000100111011101110111011101100100011101110001011101110010001100010111001101110000011001110111001101110110011100010111001101100111001001110111001101110000000101110010011101100111000101110111011101110111011100100111011100010111010101110111011101110111011001100111010100010100000001110111011101110011011101000111001001010010000100100100000101110111011101110111011100010011001100010110000101110011011100010001001001110111001000100110",
		"01110111011101110111010001110111011100100100000101110001011101110001011101110111011100010111001000110010011101110111010101110111011101110111011101110110010101110111011101110111001001110010011101010011011101110111011101000111010100110111011101010111011101110000011101110101011101010111011101110011011101100111000001100111011101110111011101110000000001110010011101100111011101110111011100110111010001110101011101100111010101110001011001110111011100000100011101110111011100100000011101110011011101110101000101110110",
		"01010111011101110101011000010000010001110111011101110110001101110111001101110001011101110011011101100111010100000111011101110010001001110111011101010101011101110111001101100111011000100111011101110001001001110110010001110111011001110110011101110111011101110111011100000110011100100101000001110111011101110111011101110111011100010100011101110111011101110111011001110111000100100111010101110111011100000111010001100101011101110111001100110011000001110011011101110000011101100100010001110111000101110111011101000011",
		"01110001011001000111011101110111011101110111010101110111011101110111011100000011011101110000011101110111011101110100011101110110011101110001001100010111011100100111001101110000011101110000011101110111011101110111011001100110011100100111011100110110001101110011011101110011010100000111011001100111011101110100010001110100000001110111000101110111011101010111000101110101011101110100000101110111011101110001011101100111011101000011011101110111010000000111011101110111011101110111011001110111011101000111011100100111",
		"01110010011101110010011100110111011101110101010001110111001101110000010101110111010001110010000101110111001101000111011100100111011101110111010001110111011101100111011101110001011101110110011101000111011101110001011101110111011001000111001101110111011101110110011001110110011100000111011101110111001001100111011101000111000100010111011101110111000100000100011101100011000001110111000001100110010101110111010100010101000101110011011100000000011100100111011101100100011101110111011101100111001001110000011100100111",
		"01000110011101100111001001110111000101110111011101110111011101100110000101010110011001110101011100010111011101110101011101110111011101110110011101110111011100100111011101110010011101110101011101100111011101110111010100010111001001110111011101110111000101110010011100000111011101110100011101110010001101110111011101110011011101110001011100010111011101110111011101110110001101110111011001100111011101110100000001110111001000010011011101110111011100010111011101110010011000110111011101110000000001110011011101110111",
		"01110111010101110111010100010111001000000010011100100111011100110110010001110111011101110111000000110011011101110110010001000000000101110111010101110111011001110111001000110111011000100100001001110111000101100100011101110100001001110000011101010111011101110111011101110110000101110111000001110111011101110110011101000111011100100111000101100111011101000110011100010010011000100000011101110001011101110010011101110111011100000001011100100111011100010001011101110111011101110011001101100111011101110011011101000111",
		"00010111011100010111011101000111011001110100011101110100011101000111011101110111011101110001011101110101011100010001011101110111011101110000011101000111011101010010011101110111011101110101001001110001011101110111011101010100000001000100011101110001011100100111011101110111011101110111011101110111001101000100011101110111011101000111011101110111011101110111000100110111011101010111011101110111011101110101010001110111011100000011001101110111010001110111011101100101011101110111011100000111000101010110011100000111",
		"01110101000000110111011101110101011100110110010001110111011101110111011101110111011101100111000101110111011101000010000001110111000001110110011100010010011101110111011001000000011101110101011101110111011101110111011101110111011100110111000001110111011101110111011101100101010101110010011100000100011101110111011101010111000101110111011101110111011000100111011100000111000000000010011101110111011101110111011101100000011101110111011001110111011101110101011100000010000000100111011101110010011101110111011101010111",
		"01000111011101110001011101110111010001110111010100110111011101110111001001000111011000000111011101100110011000100101011001110000011101110111000101110000011000010111000001110111010100000111011101000111000001110010000101110010011101110011000000110000011101110101011101110111001000000100011100100111011100100111011101110001011101110111011000100111000000010111011100000111011100100100011101110101011101000111011101010111011000010011011101110010001101110111011101110111011101110101011101110001010001110111000001110001",
		"01110111011101110111001101110010011101110100011100110111000001110111011001110110011001110111000000100011000101110100010001110111011100100110011100010100011101110010010101110111000001110111001000110111001000110111011101110001011101110111011101110111011101000001001000100010001101010111011101110111010001110111011101110111000100010001011101110111011101110100000001110111001001110111000001110011011001110100011100010111011101010111011101110111001101010111010101110111011101010010000101110010011101010101011101110111",
		"01110111011101110111010101110111011101100111000101110111011100110101011101000111000100000111000101100111010101110111011101110111011101110111000001110111011101100011011100000101000001110111011101110010011101010111011101110111011001110111011101110101011101110111011100100101001101110111000101110111011101010010001100010010011101110101011100000111001001100110001001010111001001110111011100100111011100100111000001110111011101110111011100000011011101110100011101110111001101110111010000110011011101110001001100000111",
		"01110010010001100010011100100111001101110110011101110111011101010111010100100111010001000111001101110010011101110111011100000111010101010111001101110111011101110111011100000110010101010011001100100111011100110111011101110110011101110111011101110111001000010111011100000111000001000000011100010111011100100110011101000111000000100111011101110100011100100011010101110111011101110111001101100111010000100111000100000110000001110001011101110111011001110101011101110111011101110111011101010001011101110001000101010111",
		"01110111011101110111011100110001011101110111001101110111011101110110010101000010000101110111011101000111001001110010010000000111011101110111010000000100001001100011011101110110011101110111000001110000011101110110001100000111011101110101011101110010001001110111011101100111011101010111010100110010011100110010010001110111011101110111011001010010001100100011010001110111011101000100011101110111001001110111011100000111011101110101011101110111001001110111011101110111011100100111011100100101000001110111010001110111",
		"00010111001100110000001001110001010000000111011100010111011100000100011101110111011101110111011101110101001001110111011101110111001001100000010001110111011100000111010000110101001000100111011101110110011100010111010100110111011100110111011101010111011100010111011101110111011101110111011101110111011100100011011101110011011100100011011101000111011101000100011101110111011101110111011100110111011101110011011101110111011101110011011001000010011100110111011001110111000001110111011001100010011101110010010101010010",
		"00110111011101110111011001110111011101110111001101000111011101110111011101110100010101110111010001110111010001010111010101000111011100100110010101000111001001110111010101110111011100010100011100100111000000110010011000100111011101110111011100000111000100100111001101100111011101000000011101010111011001110111011001000010011101010111011101110011011100110101011101110111011101110011010000100010011101110111011001110100011101110111011101110101001001110111011100000111010100000111011101110111000001000010011101110101",
		"01010111011100000011001101110101001101010101011001110111011101110111011100110110010100010001000101110111000101110111001101110000000001110111000001110101011100110100011100110100011100110111011100010110011101010110000101110111000101110111011101110111011101000111011100000000011100000111011101110001011101110001011101110111011101110111010101110111011100010010011101110011010000100111011101000010011101110101010001100011000000110011000000000111011101100110001101010001000100000111000101110011011100110011011000000010",
		"01110111011101110010011101110111010101110111011101110111001100100001011101110111011101110001011101110111010001010111011100000111000100100110011101110001011001010101000101010101010101000101000101110110001000110111011101110111011001100111011101110111011101110111011101000100001100100000011101110111001101110000000001000111011101110000011100100010011101110110011101110111001001110111011001110111001000000011010001100111000100110111011101010111011101110111000101110111011101110111010001110111010000010111001101110001",
		"01110001011101110111010001110111011101110111001101110111010001100111011100110101011101100111011101110111011101110111001000010111000101110101011101110100000001110101000001110001001001110011011100000111011101010111011001010111000001110001001101110111011101110100001001110111011101110111010001110110011100110011011100110100000101000001011001010000011101110000011100000111011101110111000000000001010100100111000001110111011101110111011000100110011101110010001101110111011101110111011101110101011101110111011100110110",
		"00100010011001110011011101110111000001100111001001110010011001110111010101110001000001010111011001110111011001110001011101010111011101110111000100100000011101110111000100110000011101110000011101110111011101110000001000100111011101110111011101110111000101110111011101110111011101110100011101110110011001110111000101000010011100010111011101110111011101000111011101110111011101110111001101110101011101110111011101110101011100110101011100000010011101110111011101110101011101110111001101110111011101110111010001000111",
		"01110111001000100001011000110000011101010110011101110111011101000011001001110111011100000010011101010111011101110000011101000111000000100111011101100111011101110111011101110111010000000111011100010001011101110111011101110111010100110111011100000011010001110111000001110100011100100111011101110111011101110000010000010111011100110111011001110101011100110111011101110111011101110110001101110111011101110111011101100111011101110111011101010111010001000101011101110111011100010111001001010111000001110100001001100111",
		"01110111011101000111011101000111011100000111011101110111011101110000011101110011000101110111011101000111010100100111011101110111011001110111000101110000011101010101010101100111010100010100011100100001010101110111011101110000011100110000001001110111011101110010001000110111000101110111011101100000011101010111001100110111000001110110001101000111011101100111011101000111010101110111010001010101011101110111010001010111011101100111011100000111011001110111011001110111001001110010011101110000011001100100011101110111",
		"01110110010000110111000001000111011101000111010001110101011100010111010101110101011101110111010101110100011001110111011101100111011101110101011101110001011101010010001001110110011100010111010001100111011101000111010000110111000001110101011101110111011101110111001001110111011101110111001101110111010001000110011100100001001100000111000001110101000101110111010001110111011101110111010000110111011101000111010101110111011100000011011101110100011101110111001101110111011101110110011101110111001101000111011101000110",
		"00100111011101100000010001110111001101110011010100100111001101110111011001110110011100010111010000110111001101110010010101000111000100110111011101110111010101010100011100110111000101110111011101110000011101110110010001110000010101110100010000010111011101010110000000100111011101000111010001110011010001010101011001110001011101110111000101110110011101110111011101110111011101100100000100010111001101110010011101110110000001110101011100000101011101110100000000100111011101100111011101110001001101000001011100100110",
		"01110111011101110000011100010111011000000111011101110111010000010111011101100001011100110010011101110111011101110101011101110111011000110111010001110111010000110111000101100111011001110111011101110111001100110111011101110101011101110101011100000111000001010001011101110111011001110111011100100000011001110111011101110111011101110111010101000111001000100111011101110010011101000000000100000101000101110011000101110010000101110100011101010111001101110111000100100111011101110111010100110111011101110101011101110011",
		"01110111001001110110010001110111011101110100001101000111011101110000011101110100011100010100011100110110011101110111011101110101001101010100001101000000010001000101011101010101011101110000010101110111011100110111000101010001001100110001011101110111001101110010011100000101000100110111011101110101011101110111001000100011010101000010001001100001010101110111011101010111011101100110011000000111011101110110001101110101010001110110011101110111010001110111011101110111011100000011011101110100011101110111010101000111",
		"01110111000000010111000101000000011100000111011101110110011101110010010001010100001001000111011101110101011101110011011100000111010101010010011101110111011101110101011100110111011101110000011101110111001101110111011100100100011101110000011000000111011101110011011000110111011100010111001001010000011101110011011101110000011100000001011101110111011101010111011100010111011101110111001000110111001001110111000001000111011100000110011101110111011101110111000101110111011101000001011101000111010101110111011101110111",
		"01110111000101100111011001110111011100100000000001110100011101100111011001110101011001010001011101110111010100010010011100100111011101000111000001110111011101110111011100110110001001110011011101110100000101110111011101110000011001100101011101110111001001010111010101100111001101110101011100000010001101000111000101110111001101110100011101110000000001100000011100110111011101110001011100110001010001110111011001110101011100010010011101110111011101110111011101110011011101110111011000100000010000010011010100010000",
		"01110111000101110001011101110101011101000111011101110100000101010111001101110010011100010111011101110111011101110111011100110000010101000110011101100111011101110111001001110101011101110111010001110011011101110001000101110100001001110111011101110111011101110111010101110111011101110111010000000100011101010001011101110100011000110111011101110110011101010111001101000111011101110000011101110110011101110101010001110111011101110111011101110111011101110111011101110101011101110111011101110111000001110111011101100100",
		"01110001000100100101011101110100011101110111011101110111011101010111001001110000011101110111001101110010011001000001001100000100011101110111000001110001011101110111001000000111011100010111011101110111001000100111011101110111000101110001000001110111011001110010001001110110011100010111001101110111011001110111011101110111011101110101010001100111011001010111011101000001001000100000011101110001011001100011010100110110011101110011011100100111010100110111011100110111000101110111010001100111011101110110000001000110",
		"01110111011101000110011100010111011101110111011101110111011101110111010000100111011101110000000100010111000001110101011101110111011101000010011101110111011101110111011100100111001101110111011101110111010001110101011101110011000001110111011101010111011101000011011101010110011101010111010101110111011100110111011101110110010101110100000001110000011101000111011101110111011100010001010101110111000001110110011101010111001001110110001101110111010001110011010001110111000000010111000101110111011101110001001000000111",
		"00010001011101110111011101110111011101110111011101000000001001010010011101110111001000000111011101110000000100010111000001100001011100100101010100100110001101110011011101000111011100000111011101010111011101110110011101110111001101110111010001110111001001110000000001010111011100000111011100000100001100000111011101110101011101110111000101010001011101000111011101110000011101110100011101110111011101110100011100100111011101110111011101110111011100100010010101110110011101110110000100000111011101110111010101110111",
		"00000001001101110110011001110111011100010111001001110111011101110110000101100111011101110111010001010111010001100111011001110111011101110111011101010111011101110001011101110101011101110000011101010111011001110111001001110110011101110111011001110001011101110010000001110101011100110111000100000111000101110111001101110111010001110100001001110111011101000110011101110110011101110111011101110111011101110111011101110111001001110011011101110111010001110111000101110111011101010111011100000101011100100111001001100000",
		"01100111010000110111010101110111011101000110011101000000010001110111000001100111011100110100011101110011001101110111000000110011010001110111011101110111011001110111011101110111011101000100010101110111011101000111000101110011001000000111011100110111011101100010001001100111011001110101000100110111011101110100001101110111011101110100000100010111010100010111011100100111001100100111011100110111011100100111011100010111011101000101011101110111011101100000000001110001001001000111011100100101011101110011001101110111",
		"01110111011001110011011101110100011101110000011101110111011001110111011101110100000001000100001001110111011001110111010101100111011101110110011101110010011100000110011100010111010001110010011101100000011101000001011100010111011001110011010001110000001101110111011000010111011101110111011101000101011101110111011100010001010101110101011101110111001100010110011101110111011001110000010101100011001001010111011001110111010101110111011101110111011101110111011000110001011000000010001100110101010000010110011101000010",
		"01110000011101110111011101100110010001000000001101110110000001110111011101110000011101100111011100010111011100010111001101110111011101110111011101110111011101010111011100100111000101000110011100000111000001000111011101110111011101110111011101110100001000010111011101110111011101110110011101110111011100110010011101110111011100000011001000000111001100010111001101110111000101110111011101110111011100110010000001000101011101110000000101110111011100110110011001110111001101110111010001110111011101010010011101010111",
		"00000111011101110111011001110111010100000001011100010011011101110000011101010100011101000100000100010010011101100110011101110111010100000111011101110111001001110101011101000111011101110111000101100111000001110010011101110001001101110111011100110111010101110011011100000111001000100101011101110011011100010111011101110111010001110000011101110001010001000111001101110011000001110111000001110111010001110100011101110111011100010100011101110010010101110111011101000111011101010111011101110100000101110111001101110111",
		"01000111011101110111001101000111010001110111011001110001000101110110000100110001011101000111011101110000011101110111001001000111011001110111011101100000011101110111011101000101011101110000010001110110011101110110011101100111000101010111011001110110010101110111011101010111001001110111011101000000011101100001001001110011000001100111010001110101010001010010011101110010000001100111011100010111011001010111011101110111000101110111001100000000011100010111011101110111001101110100000101110111001101110110011101100111",
		"01110101011101110111001001110010001101110001011101110111011101110111011100010100011101100010011100000110011101110000010101010100011101010111011101110111000101110011010100110111011101010111001101110001001100110111011101110001000000100111001101110111011101110011001001110000011100110011010000100111011101110111011101110111001001110111001101100111011100000111011101110100011101110010011101100001011101010111000000110111010001110111011101010111011101110010001000010111010001110010011101000111011101110111011100000111",
		"01010111011101110110010001110110011101110111000100100111000100100001011100010111011000100110011101110010011101110111001101110111011101110111011100010000010100000101011101010111001101110001011101100111011100000111011101000111011101110001011101110110011100000110011100110111011101010111011000010010011101110111000001110111010101110010011101110011011101110001000101110111011101100000000101110000001101110111011101110111011101110000011101110111011100110111001101110111010000110111000001110111010001110111011101110110",
		"01110111011101110111010000100111011100100100011101110111011001110100011101100100010001110111011100100111011100000000011001110111010000010111000001110111001101010111011100100011011101110101011001110111011101110111001001110111011101000111011100000011000001110111011001110101011101110111001001100111011100000111011101110110000101010111011101110111000000100100011101110111000001110000011101110100010101110111011101110100011001000011011101100111011101110100011101110111010100110111011001110110010001110101011101110111",
		"00010111011100110100000000010110001001100111010101110011010001010010010001110101011101110110001001110111011101010101011101100111011101110001011101110110011100110111000001110111011100100100011100110100011101110101000101100111001001010000011101010001000001110010001101110111011101110000011001110000000101110000010001110100011101100111011101110111010100010100011101010001001001110111011101110111011101110010011000110000011101110111001101100001000101000111001101110001011100010000000101110011011100110110001101110001",
		"00110001011101110111010001010000010101110101000001110111011100110110001101110111011101110111011101110111001001110111011101110111011101110000000100100111000001000011011101110010001101110101011101110111011101010001011101000110001001110111011101110111011101010010011100010110000101110111011100000101011101110111011101110001010101110001011101110001011100100111011101110111011101110011011100110011010101110001011101110010011001110111010101010010011100000100011101100101011101110001011100110011011001110111011100110110",
		"01110110010001010111011100110111000001110111011101000101011101110111011101110111001001110011001001110111011101010010011101110000011101010000000000010100010101110111010101000001001001110111011101110000011000010011001001110001011101110101011101110100011100110111011101110111011101010000011100110100000001110111011101110111011101110111011101110111010001110110011101110001011100010111000101110010011101110111011101110111001101110111001001000111011101110111011100000111011101110111011100100100011101110111001101110101",
		"00110111011101110101011100010011010000100111000001110110011101010100011101110111011101110111001101110010000001110111011100100101011101110100011101110000010000110111001101110101011100000111000001000111011101110111011101100111011101110010010101110010011101110101010000000011011001110111011101110111011101000100011001110111000101010111011101110011011101110111011101110111010001110111011101110111011101110110001001110111011101110111011101110110001101010000010001110111011101110011000001110111011101110100000101000100",
		"01110000001000000001011101110010001001110100011000110111011101110111000000010111000101010100011101110001011101110101011101110111010101110111000001110111011101110011011101110111000001100100001001010011011101110111011100100011011101100111011101110011011101110111010000000111000101100111011100100001011101110111011101110001011001110111011101110000001101110000011101000111011001010111011101110111011101110111011100010100011101110111001001110111011001010111011101110111011101110111011100100111010101110111001101110111",
		"01110111010001010000011101110001001101110111011100100010011101110111001001110100011000000000010001110101000001010111000001110111001101110111011101110100011100010111011101110111011100110101011101110100011101110111011101110100011101110100011101110111011101110111000100110111011101000000001000110100011101110010011100110000011101110111000000110111001001110111011101110111011100000111011101110111011101110101001101110111011101000101011101110001001000000111011100110111000101010110000100100111011101110111011101110111",
		"01110111011101110011011101100111011101100111011001110000011101110011001101110111000101110111011101110111001001110100011001100111011101110001010100000111011101110111011101110000011101100000001101110111011101110111011101000111010001110111011101110111011101010111011100010111000101110111001101110010000001110001001000110010011101110111011100100000000100010111011001110111011101110010011101110010011101110111000101110111001101110111010001110110010100010111000100000111011101110111000100110111011101110111000101110111",
		"01110111000100110111011101110111011000100111011101110111010101110111011101110111011001110110011100110111011000000111010101010001011101000111000001110111011101110000011101110111011101110111011101110111010101110110011101110110010000110011000001110001011100010111011100100111010101110111000000100101011100110111010001110111011101100111001100100010001001010011001001110111011100110111010001110011011101100111011101110111011000010011011101110000011100010010011101110100001101110111000001110100011101110010011000010111",
		"01110111011101110111011101110111011101100010011101000110011101000001001001010101011101110111000101110011011101110010011101110111011101110111011101100111011000110111011101110111011100100010011101110100011101010111011100110111010100000101000101110111010000000111010101110100010101110111011100100111011001100111001001110101010000110101010001000110001001100111011101100110011000110111010101110111000101110111010101110111011101110111010001110011010001100001010001110111011001110111011101100111011100000111001101110111",
		"01110111011101110111010001110110000001110110011101110111011101110010011101110111011001010110011101110110011100000010011101110100010101110100001100110011011101110111001101110011011101110111011101110111011101010001011100010111000101110110000000010010011101110110010001100111001101110001001101110010011101110111011000110001000100100111001001110110011101110000011101110110011101110110001000100111000101000100011100000111011001110111011100110001011101110001011101110111010001110101010001110111000001110111011101000010",
		"01110001011101110111011100100111011001110111011101110111011101110110000101010000011100000001011001110011011000000111011100010000011100010010001101110110011101110111011101110111011101110111011101110100010000110111000001110010011101110001011101010010011101110111000001100111010001010111011101010111011101110001000001000111011100000111001001110111000100000011001101010111011100110010010001110111010101110100011100110111000101100111010000100111011100100111000101110111010001110001000101110111011000110110011101110111",
		"01100010010101100111001101110111011101010011011101110111011101110101011100010111001100100111011100100010011100010000001000000111011001110111011101110111011101010111011100100111011101110111011001110111011101010000011101110100000000100010000101110111011101110111011101110011000000100111011101100111010101110001011100000001001001110101011101000111011101110110011101100001011101110100011101110111000101100011011101110011001001000111000101110111010001110100011100110110010101100111010101000100011001110010001001110001",
		"01110110010001110111011100110101011101000111001001010111011101110111011101000000011001110111011101110111011100110101010101110110011100110111011000110111011101110111011000110111011101110111011100110111011101010111010001110011010100110111011101110111011101110111011101110111011101110111000101110111011101110100011101110110011100100111011001010001011101110111011100100111011100110111001000000110011101010111011101110001011101110010000000010111010101110010011101100010011101010011010101000100001100000111011101110000",
		"01110111010101110001010101110110011100000000010001100111001101110111011100010111011100000100011101110111011101110111010001110100000001100111010100110000000100110110011100010100011100000010011101100111000101110101000101110000001000010000001001110000011101110111011100100101011001110001011101110111000000010101011101110111011101010111011101110111011101100111000001110111011100000111011100010111011101100111000101110111001001110111011000010111010100110111000100110010011101110000011100100000011101110111011100000111",
		"00100111001001110111011101110110011101110010001101110010011100100101010100000111000101100110011100010011011101110000011101110000011101110111011100110110011101110001010000000111011101110001011000000111011100100111010100000111011101110001001000010101011101110011011101110111000101110111011101100111011101110110011101000111001001110011011101010111011001100100011101110000010101110111011101010111011101110111001001110101000100010010011101100111011101100111001001110111001001110111011101110111011101110010000101110101",
		"01110101011101100111011101010000001001110011000100010111001101100101011101100111001101110111010101110110011101000111011101010111011100100100010100100111011101010111010101110111001001110000010101110111000001110010011101100111010001000111011101110111011101100010011100010111011101110111011101110101011101100100001001110000011101110000011101010111010101110111011100110111011101110110011100010111011101110111011100000111001001110111011101110000011101110000011100010001011101110101011100100101011100000111011101110111",
		"00100111011100010111001001110111011101100111011101110111010001110000011100010010011101110111011100110001011101110111011101100111011100100111010000000110011101110111011101110111000101110111011001010011011101110111011101100101001001100111011101110101000000000101010101110111011101110111011001110010011101110110001001110001011101110101001001110101011100110111010001110111000101110110000001110111011101110111011100100011011101100111010101110111011100000111011101110111011101110111011101110111011000100101011101110111",
		"01110111011101110000000100110011011101110101011101100111010100010111010001110111011100100100010001110110010000110111011101110100011101110111010000110010011100000111011100100110001001110111010101110111011101100101000101110111011101110111011100110111011101110111010001010111011101110001011100000011011101010110011101110111011101110111011101110011000101110111011001110111011101110111011101110111011101110111001000010111011101110111011101110100010100010111010101000111011001110100001100110111011101110111011100000100",
		"00010001001101000010000100000000011101010111011100100111011101110111011101000111010101110111001100110111011000010011011101110111010101110011010101010000011101110000011101010011011101000111011101100111000101110111011100100000010001000110001101110000001101110111011101110011011101110010011100000111010101110011011100000001010100010111011101110111010001110110011101100111011101110111001001110111010101110011001001110111011100110010011100000100011101110101011100010000010101110111001001110111010001110111011100010110",
		"00110111011101110111011101110001011100010111000101110111010101100110011101110111011100100111011101110000000101110111001100100111001101110100010001110010011100000111011101110111011100110111011100110110011101110101011101110110011101110111000101110111011001110111011101110111011101110011011100000100011101100111011101000111011101110011011101100111011101010101011101110101010101110110011101110011011101110111011101110111011101110111011101010110001101110111011100110110011101110111011101110110011100110101010000100111",
		"01110001011101110111010101100111010001110111001101110101011101010111010101110111001101110111011101110100010001110100011101100101011101110100000101110001010001110111011101110111011100010111010100010111011001110101010101110001011100000110011101000010011000010111011101110010011101110111001100110110011100000111011101110111011101110011011101110100001101100000011101110111001001110100011101110111001101110011011100010111011101110111011101110011001101110111011101100010001001000100001101110111011001110111011100110100",
		"01110111011100000111011101110101011001110110011100110000010101110000001001110100011101110000000101110111001101110000011100010111010101110001010001110100011100100111011101110010001100100101000100010011011101110110011100100111011101110111011101110111011101110111010001110101000101110110011101110111001101110111011001100111010100100011011101110011011101100001011101110111011101010111011101110001011101110111010100110111011101110111001000110110011101110111011101110111011001110111011101110111000100000101010001110010",
		"01110100011101110111011001110111010101110111001001000111000101110011011101110111000001110111010001110111000001110111001000010111011101010111011101100111001001110111011101010111001101110001011101110111000000100111000101000101011101110111011101000100011101110111011100110111011101110111010000110111011101100111011101110111001001110111011101110111000000010111011101110110000101110111000001110111000000010111010001110111011101000111011001110101010001110111011101000001011100010101010000000111011101000000011101110000",
		"00000111010001110100001101010111000101110101011101110001010001110110000100100001011101110111000101110111011101110100000101100101011000000111011101110111011101110111011101110111010001100110011101110101011101110111011101110110001101110110011101110111011101110110000101100111011101110011011101110111011101110111011101110010010101100111011101110011011101110100011100010101000101000100011101100111011101110000011100110111000001110001011101110111011101110010011101110010011101110000000001010011010001110101011001000110",
		"01110010011101110111011101110111011101110111000001110111001001110111001100100111011101000111000001110010011101110010011101110111011101110000000001110111011101110000011001110100000101110010011101010111011100000111010001000111000101010100011101100111011101110111010101110111010001110010010001110100011101110000010001110111011001100110011101100111011100000111011000010111001001110111011100100111011101000111011101110111011100100111011101110111011101100011000001110111011101100000000000110111001101110111011101110111",
		"01110101011100100111011101110000011101110101001100110110011100000100011100100111011101110111011101110111010101110111011101110001010000010111011101110010011101110111011101110111011101110111011101010111000100100010011100010100011101110001011101010000011100000100001000110111011101110111011101110111011101010110011101110001011101110111011101000011000101110111001000010011011101110010011101110111011001110111011101110111011101110111010101110011011101110111011101110111011101110001010101110111000001110111001001110010",
		"01110111011100010111011101110111011101010111011101110111010101110111001101110011010001110111011101110111010100100010011101110111011100000111000001110011011100000111011101110110010001110111011101110100000001110111000101110111001000010101011100010111011101110000001001110110000101110110010101100000011101110111011001110111011101110000011101110111011101110110011001000000011000110111011101100111001101110111011100000000011101100100000000110110000001110111000000100111011100010011011101110010000101110111010101100111",
		"01110011011101110010011101110111010101110011001101110111011101110111011101010111011101110111011100110111011101110111010101110111001001110111011100000111011101110110011101010111011101110111011101110111011101110111011101110010010100010111011101110101000001110010011101000101000000000111001100110000011101110000011101000111000101100011011100100111011100110111011101000110011101000011010101000111011101100011010000010110011101110111011100000111010101110110011100100111011100010111011101110111010100110100011101010111",
		"01110111011100100000010001110011010100110111001000100110000001110000011101110111011001010011010001110111010001100100011101110111000101100111011101100111011100000110001100000000011101010110001101110111011101110111011101110111011101110111011101110000011001110111000001000111011101110001001100100111011100110011011101010111011000010001000001110111000000000111011101110111000001110111011101100111011101110111001001110111011001100111011100010100011101110110001001000111011100110111011100100010011101110111011001010111",
		"01110111001101110111010101000001011100000101000001110111001101110111011101110111011101110111000000110111000001110011010100010101011101110111011100100010010101110111000100010110000001110001001001110010010001110011000001110110001001110111011101110111011101110110011100010111000001110000011101110100011101010011011100000110011101110000001001110110011101010000001101010111011000110000011101110111000101010111011101110111011101110011010001110111011101110111011101110111000001110001000100000100011100010110000001110011",
		"01000111011101110011011101110111011101100011010000000111010001100111011100100111001001100001011101010111001100000000011101110111010101110101000101110010000000100010000101110110011100100110011101110111011100010111011101110111000101110111011101110111011101110111011101110010011100110010001101100111000101110111011101110011000101110101011101000111011100000000011101110001011101000011011101110111011101100000011101110010001001100111011101010100011101100111011101010111001100010110011101110100000101110001011101110111",
		"00010111011101110111011101010011011101000111010101110111000001100111011100000111011101110001011101110111000001110011001100110001011001110111011101110001000001110111010000000111011101110110011000110111000001110000011001110111011101100100011100010111011101110111011101010010011101000000011101110111011101110010011101110111010100000000011101110101011100100111011100000101011001110111001101110111011100000111010001110111001101110111011101010111001101110111011101110000011100100111010001110111011101110011011100110111",
		"01110111010100000111011101000111000000010111000100000100011101100111011100010111000000110111011100000111011101000001011001110111000001010110011100010000001001110011011100010111011101000000011101110110010001110111000001110110011101000111000001110111011101010111000000110111011001100111001101010111011100000111011101110111000100100101011100110111000101000111011101100011011101110111011001110111001100000111011101110010000101110111000000000111001000000010011101000111001101110101011100010110001001110111010101110111",
		"01110111011100110110011100010111001001110111000001110011000001110111011001010011000101100111011101110111010001110111011100110111011101110111011100110100000101110000011101110110011101100111001100010010000001110000010101010111010100100111001101110111011100000110001101110111011101110111000001110111011100110100011001110111011100100111000101110011011100000010001101110100011100100001011101110100000001110110011101110001011101000010011100000001011101000111011100110111011100010101011100000000011101110111011001110000",
		"01110111010001110001011101110011001001110111011101110111011101110000011101110000011101110110011101110110001001000111011001110111010101110111011100010101001001110111000000110111011000000010011101110000011100010101011000010111011101110100011101110110010101110000011101110111001001110011011100100111011101110011001001110111000101110000011101110111011101100111001000010111010001110111011101110111010001110111001000100010010100010011011100100111011001010111000101110000001100110110011001000111011001110101000101000111",
		"01110111011100000111011101110111010000100100011100010100011100000101001101110111011101110111010101110111001100010111011101110111010001110111010101010111011101110011011001010000000001110111011101010010001000110111011101110111011100000110011101110111011101110111011101100111011101110111011101110111011100110001011101110111011101110110011101110111011100000010011101110100010000100110011001110101011100110010011101110111001001110111001101110100011101000111011101110111011100000011011101110001011101110111011101110000",
		"00010111011101110111011101010111010001110111011101110111001001110110011100100111010101110011011101110100011100100111010000100111011101010101011100000111011101110110011101110111011100110111001001110111011101110101011101110011011000000111011100110110010101110111000101000111011101110111011001110111011100110111011101110111011100100001001100100111011101110101001100000111001101110111000100110111011101110111010001110111011101000010011001000110010101110100001001100111011101110111011101110011011101010010011101000111",
		"01110000000101110111011101110111011001110111011100110111011101010111001001110110011101110110000000110111000000110111011100100111011101110011011101110111010001110111011101110111011101110111000001110111000101110000001000100011001101110111001001110111001001010111001001110111011001110111010101110111011101010111011101110111011101110111011101110111001000010111011101110111011100110111011100000111011101110000010101110111000001110101000000010111011101110111001000100000000001100111000000010110010101100000011101110110",
		"00000011011101110011011101110100011101010111001101110111011101100110011101110101011101110011011101110111010001110010011101110111011101110111011101000011011001110110000000010111011100100110011101010001001101110111011101110100011101110111011101110111011101110010000001110111011001110111001001110110011101010010010101100111011100010111011101110110011101110001011100100111011101110111011101110111010101110111011101000111011101110111001101000100010001100111011101110111011101110010011101110000011101110100001000100111",
		"00010111011101110010011101010110011000100010011100110111011001110000011100010111010001100101001000010111011101110111011101110110001100000111011101000011011101110001011100110111011101000111011100010001011101110000011101110111011101110111011101110111011101110111011100100111010101100111001000110111000101110111011101110111011001110111000000010011011100110101011100110111010001110011011100100100011101100100011100100101011100110100011101110111011101110100011101110011011101110111011101110111011100100111011100000111",
		"00010011011001110001000001110111011101110111010001110111011101110100001000010111011101110011001100100011010001110111011101110111011101100111011101110111001000010101011101110111010001010001011100000011011101110000011101110111001101110001011101000111011101100100011101000111011100000111011101110111011100010111010101110110011101010101010101010111011100100111011101110111001001110111001101000011010001110111011101110001011101110111000101110000011101110000010101000111011101110111010000100001011101100111011101110101",
		"01110111001001110111011101110111010001110111010100010101010101110000000000100010011000010010011100010111000101110111011101110010011101110011011101110111011001110001011001110111000001110011011100000111011100000101011101110100011100110100000101000111010000100100011001110111010001110111011101110111011101000111011101100111011101010110011101110001011101110111011101110110011100110000011101110111011100110111011101110111011100000111011100100111010101110111010101100100011100110111011101110111001100010011011101010001",
		"01110001011100110010011101110111011100000001011101110111011101000101011101110111011100110111011100010111001001100011011001110001011101100111001001100111010100000111011001110111011100110010010001110111011101110001011100000010011101110111011101110111000101110111010001110111001100100111010001110111010101110000001100100110011100100111001100100111011101010011000001110011001000100011000001110111011101110101011101110110011101110011011101110111011101110111000001100111011101110101011101110001011101110100011101110111",
		"01000111011101010001011100000110010101110100010101110111010000010111011101110010011101110111000101100011011101110111011101110000011101100111011101110111010101110111011100000010011100100111011001000111011100010111011101100111011101110100011101100111011101010110010000110110011101110101000100100111001101110111011000000111011101110000010001110001011100000110011101110111000101110100011101110111011001110010011101110111011101110111011101110011011101110011011101110111011100100101000101110111011101010111011100010111",
		"01100111010101110111001001110111011101110001011101110111011101110111010101110000011101010001011001010111011100100001011101110111011101110100001101110111011101110111011101110111011000100111001101110100000100100110011101100001011101110100010001100111011101010110011101110100000101110100011101010111011100000111011101000111010001010110011101110111001101110000001101110100000001110111011101000111011101110000000101100111011101110100001100110010010001010111000001110111000101110001011101110111011001110111010000110111",
		"01100011011100010111011001100101000101110110001101110111010000110101011101110000000000110011011100010111011101110101011101110111011101110011001001110111011101110111000101110000010001110111010001110010001001000111010101100111011100000111000101110111010001110111011101110101011101110010001101100111001101110100011101010111011100000100001101110010010100000111001101110011011101000111011101100101011101110101001101110111011101110110011100010000011101010100011101110111000101110110011100000111011101110010001001110100",
		"01110001000001110111011100000111011101110100001101110111011000100111011101110111000001110010011000000111000000100100011101000011011001110111000100110010000101100111011100110111001100100111001101000011000100110111011101110100011100000111011001100111010001110111001101110101011100000001001001110011010100010111001001000111011101110101011100010111011000010100010101110111010101010000010001010110001101110100010101110111010101110011011101110010001101110111011101010111011100100111011101000111011101100111000000100111",
		"01000111010001000001000001110000010000100111000101110111011101110111011101110001010000110111000100110111011001110100001101110111001000110111011101110111011101000111011101110111001101110111011101110000011101110111010101110100000101110111011101110111011101010010000001110111011100110001011001110011011101100111011101100111010101110100000000110111011100110111011101110111000101110001011101110010011101110010011101000111011000110111000100000111011101110100001101110111011101110011011001000111011101110111011101110010",
		"01010111010101110111011101110000000001100111011101110111011000000111001001110111001101110111011101100111010101110111010001110111001001110111010001110001011101010100001001110111011101110111000001110111011101110101011101110111010001110111000001110010011101010111010001110001011101110111000100110000011101110001011101100111001101110010011101110111001001110111001101010111011101110111001101010011011100100000011100100111011100100000000101110011011100100110010001110111011101110001011001110000011101100111010001110111",
		"00000001011101110111010101110101001100010111011001110111000101110111011101010111000101110111011100010101011101010111011100100111011101110000011101110000010001000111011101110111011001110111001001110100001100010110000001110111011101110111011101110100001001110111000001110101000001110111011100110111011100000111011101110111011000110111011101010111011101110111000101110001011001100000011101100111001000100010011101110111011101110111000100110011010100000111011100110111011101110010000101110111010100110111011101110111",
		"01110111001101110111001101000111011001110111011101110001000101110110001001110001011101110101011101110100011100000001011100000111000001000000011101110111001001000001011000110111011101110111011101110000000101110111011100010101001101110111011101110001011100000111011101110110000101110111010001110101000001110101001001110111000001100001011101100111010000010111011001000101011101110111001101110000010100010010011101110111001101110111011001110111011101100111000100110101011101110101011101110111000000110101011000100111",
		"01100111011101110111011101110111011101100111011101110111011101100111000001110111011100010111011101110001011101110111001101000000011101110111011101110110011101110111011101110111000001110111010000110110011100010010011101110111011101110111011001110101011101110111001001110111000001100011011101000111001101110110011000100111011101110111011101010111001000110011011101110000011101110100010100100111001001100111011101110101000100010111011101110111011101110111011101110111000001110101010001110111011101110111001101110000",
		"00000110011100000110011101110000011100100111011100110101011001110011011101110101011101110111011101000111001001110111011101110010000000110111011101010111001001110111011100010111000101110111011101110111011101010010010101110101000000010000000001100110011100110111011101100111000001110101011101100111010000010111011101110111011101110111000001110111011101110111000101110100000101110111010001110001011100110111010001010111010101100001011101100111001101110101011100100110001000000011011101110111010001110101011101110111",
		"01110111011101110001011100100011011101110111011101100010011101010111011101110111001101110000010000100010011100110111011101110111000000100111011101110111001001110111000101010100011101110000001101110111011001110001011101110111011101110111011100000111011001100101010101010111011100110000011101110111000100010001011101110111001001110111001001110101010001110001011100110111010001110000011101000010011100110111011101110111011101110000011100000111011100010001011001110001000101110110001001110010011101110111000100110111",
		"01110111010000000001000101110101011101110111011101110010011101110111011101110011011101110111010001010100000001110110011101110111000000100111011100100000011100010010011101110111011100110111011101100111011001110111011101000111011100010011011101110010011100100111011101000100011101000111010101110111011101100111011101110111011100100111001001110111010101000111001001110100010001110010000001110111011001110111011101110000010001110101001101110000011100100111001101010000011101100011010000100100001100010101011100000001",
		"00110111010000110111010000000011010101110111011100000111011101010110011101110111011101110101011101110111011100000111011101110101011101110111001001110010011101110111011101110111011101110111011101110111010101110111011101000001011101110101010101100101011101110111011101110111011001110111011101110111011100100011011101110110010001110010011101110111000100110111011101110001001101110110011101110111011101110111011101110101011001110010010000010111011101110010011101110111011101000101001001110001011101110100000100100111",
		"01110111011100000111011001110100010001100110011101110000011101110100011101110111011100010101010101110111001101110001001101110111011101000111011101010010001001110111010001110111011100000101011101110111011101100111011101110111011100100001011101110101000001110111011101110101001001000000000101110101011101110111011000010100011101100111010001110101010101100010001100100111011000000100010000100111010000110111011101110101011001110111001101110111011101100111010001110111011101110010001100010111011100010111011100100111",
		"01110001011001110101011001110010000001110100011100010111011101110111001001110110001001110111001001010101011100010001011101110111011101110111011101110011000001110111000100110111011100010101011100110101011001110111001101110100010101100101000101110000000001110111011101110100000001110111011100000111000001100011010101110111011101110111001101110111011001110010010001110111001001110111000100100110011101110001000101110111011101110111000101110111011101110110011100010111011100010000011101100011011101100111000101100000",
		"00010111011101110111011100100111010000010110000001110111000101000111011001110111011101110111000100000111011101110001011101110111010000010111011101010011011101110101011101110111011101110111001000100000011101110010001101110011011101110111000001110111011101110101001101010111000001000001010101100000000101110001000101110111011100010100011100110111011101110010000000100111011001110000011101110111011101110111010101110101000001110111011101110111001101110101001101010100011001110001001101110111011001110100011101110010",
		"01100111010101100111011101110110011100100111011100000010001000110100001001110101001000000111011101110101001001100111011101110100011101110001011101110110011101110111011100100111000000000111011101110111011101110111011100110111011100010111011101110111001101110010011000110111010001110111001001110111011101110111010101110111011100100111011101110111011101100110011101000011011101110111011101110011001101110001011101110000011101110111001000110111010101110111011101110111000001110111011101010110011100100111011101110111",
		"01110001001101010000011101100111011101110111011101110111011101000111011100110111011100010111011101110111011100000111011101110111000001110100011101100111011100100111011101110001001100110011011100110111010101110111011101110100011101110111011101110111011101110001011101110111001001110111011101110111001000010101001101110000011100110111000101100111011101010111011101110101011100100111011101100111011101000111011100000111001001110111011101110010011100000111011100100111011101110111011101100111011101110111011101110010",
		"01110110011001110101011101110100011101000111011101000100011101010101011100010001011101110111011101110001011101110111011101110110011101110111001101010010011101110101010001110000001001110101010101000001001001000111011100010111011101110111011100010111000101110111011101110110010101110000000101110011011001110111001101110111011100110010011101110100011101110101011101110111011101110111000001110111001000110001010101110100011001110111011100110101001000000101000000110001011101110111011101110111001001110111011101110101",
		"01110111011001000110011101110110000101110110011101110111011101110111001101110111010101010111000001100111000100100110011100010000000001110110011101010111000001110001011101110100001100110100001101010100000001110101000001100000000101110001011101010011011101110110011101100000011101110010011101110001011101110011011100100101001101000010001000010111000000110000011101110111011100100111011101110111001101000100011100100111011101110101000101110111000101000111010001010100011101100110010100000111011101110111011101110111",
		"00100111011100000001010001100111011101110111010100010100011001110111011101110111000001110111011101110111010001000111011100110000000101110000011001100010011101010111010001010000011001110000011101110111000101110000011100110111000001010111001101110010011000110110011101110111011101010111011100000011011101000111001101110111011001110111011101010111011101000000010101000000011101110111011101110010010100100101001101100111000001110001011100100011011100000111011100000101010101110111000000010111011100100101011100000100",
		"00110100001101110110010101110111000100010001001101010111010001100111011100000111001101110111011101110111001101110111000001110010010001110111010101110101010100000010011101110111011100110111010000010111011001110111011101110111001101110111011101110111011101110111011101110111011101110111001001010110011100000111000001110111011101000111010101110100000101110111010001110111000001110101010000000100011100110111000100000111001001110111001001010011001000000111011000100111011101110011000000000111011101000111011101100111",
		"01110111011101110010011101100111011101110111011100010000011100100110001000110111011100000111011101010111010101110111011001110001000000100111010101110011011101110111011101110111011101110111011101000111001001110111011101000111011101110111011101110010011001110111000100100011011100110011011101110101011101110111011000010111011001100100011101110101000100100111001001110111001001110011011101110101010001110111010101000001000101110111010100100111001001110111011100110111010001110101011101110111000000100111001001110111",
		"01010110011100000111011100010111011001110011011101110111011101110100011101110111010100010101010001110111010001110111011101110111011101000100011100110011001001110100011100010011011101110111011001110111011100110111011101110100011101100110011100010110001001000111010101100010011100110110011101110100011101110111011101010100011100010011000101110010011101110111011100110111010001110101011001110111011100010010011101110111001101110011011100010100000101110111010001110011001100110111011101110111011101110111001001110111",
		"01110111011100010111011101110001011100110111010100010111011101110111011101110100011101110111010101010010000100100001011101110111011101110111011101110111011101110100001001110100000000100111001101100010011101010000011101100110001001110111011101110111011101110111010001110101000100100111000100010101011100100100011101000111011101100000011001000001010101110011011101110011011101110111010100000011011101110001011101110111010001110011011101110111011000010111011100010111011001110111001101110011001100010101011001110111",
		"01010111011101110110011001110011011101110000011101110111011100100111001101110101000101000111010001110101011101110110001100000011001001110001011101100111000001000100011100010111011101110110011100110010000101110111011101110110010000000000011101110100011101100000011101110001001001110111011001110110011100110010011101110111011100010101010001110001011100110111001101010111011001110010011100000111001000000111011101110111010000100101001001110111001101110011001101000011011101110111001000010111011100010111010101110001",
		"01110011011100110100011101000111011100000111011101110111011101110001011101110111000100110111010001110100000000110001011100110101011101110111010001110111011101110001011001110000011101100111011100110111011101110111011101110010011101110000011101110111011101110111011101110111011101110100001100000011000101100010001001100111011001110110010101110111011100110111011101100011001101110101011101000111001101110111011100010111011001110000000001110111000001000111011101110111011101110111000001110111011101110100011101110111",
		"00100101001101110111001001110111010100100111011001110011001100100001010000100111011101110111001101110111011101110011011101010111011100110111011101110111011101110010011001110111011101110001011100100111011101110000010001110111011101110011011100010111010101110111000101000010011101010111001101110111011101110111000001110010011101110111011101110011011101110111011101110010000001110111010001100011011101110101011001110111000101010101011101110111011101100100011101010111000000100111001001100111011001110101010001110111",
		"01110111011101100100001101100011011101110101011101000111000001110111011101110010001100010111011001110000011100100111011101110110011101110111011101110001010100110101011100110111001000110111001100110111011101110111011101110110010100010111000101110111000101110111011101110111011101110110011101000111011101110111011101110011011101110110011101110000011100000011011101110111011100010111010001110101000001110011011001110111011101110011010001010111001100100010011101110011010101110100011101000111011101110011010001000110",
		"01110100000000000111001001110111000101110111001101100111011101110111011101110111011101110011001100100110011001110111010001110111001101110111011101110111010100010111011101110001000101110100010101000111001001110111011101110000001101110100000000110111001001110110001001110111011101010000011101110111011101110111011101110111010001110111011100010111011101110001011101110101011101010111001101100111000101110111011101110010011101010000010101110001000100110101000101110101000100100111010001110111011101110111001000100101",
		"01000010011101110011011101110111011101110111011100100011011100000111011101110101011101110001011001110000001000010111011100110111011000010101011101110111010000100111011101100000011101110101011100010111001000100111011001110010011101000111001000100111011101110111011001010111011101110111011101100011010000110000011101110011001101110100011100100100011101110111001001110100011101110111010001010111001101010110011100010111010001110111001101110111011100010100011101110111001101110011000000000111001001110110011101110010",
		"01110111011001110111001101110111011101100011011100000111011101000010011101110011011101110001011101010110000101010111011101110111011101110111011100110111011001110111000101010011011001110111010001100110011100000101011001110111000100000111011101110111011100000111000101110000010001110111011001110010000100100111001000010111010001110000001101110101000101110011011101110111011101110001001100100111000100010111011101110111011100010111001000110110011101100000000001110100011100110111001001110111011001110011001101110010",
		"01110111011101110010011101110101011100000010011101110001000000100100000101010111000101110111010001110100011101110111011101000101011101110111011101110101011101110101011101100111010100000111011101110110011101010100011101110111011101000111000100100000011100100000001001110111011100100111000001110011010101110111011101110111011101110000001001110111011100110001010101110111011101000101001001110110011101110111011001110110011100100111001101110111011101010101011101110011011100110111011101100100010001010111011100110111",
		"00000111011101110111000001110110011001110010011100000101011101110111011100110111000101110111001100010111000001010111000001110111001101000111011100100111011101110111011101110111011101110111011101110010011101110011011100010111001101000111011101000010011101110111011100110110011101100100001100000111011101010111011101110111011101110100000001110111010001110111010101110111000101100101011101110111011101110111011101110010011101110000011101110111011001100111011100010111001101110001011101100110011101100111011101110000",
		"01110111000101110110010101110110001001110111011101110011011101110000001001110110000001110010001100110111000101100011010000000111011100100100011100000111000000000111011001110111011100100111011101110111011101110111001001010111000101110010011101110111011101110101011101110111011101110100011100110111010101010000011100100100011101110111011100100011011101110101011100000111011101110010010001110000001101110111001001000111001101110111010001110100011101000001010000100001011101110111011100110111001001110111011101110111",
		"01110111000101110111011101110000010101110111001100010111011101110001011100110111011100000100011101110111011101110111011001110000000101110111011100110100001001010111011100010111001101110110000100100111011001110111000101010111010001110111011100010111011101110111010001010111011100110111011100000101011101110110011101110101011101110111001100110111011101110111011101100001001001010111011101000011011101110100010000000111011101110011011101110001011101110001011001110100011101010111000100000111011101110111001000010111",
		"01110011011101010001010101110111011101110111000100100110011101110100011101110111011101010101011101110000000101000001011101110100011001110111000100000111011101110111011101110101011101110001011101110111011101110101011100100011011001100100011101110000000101110111010001110101010101110111011101110111011101110111011001110011010001110111011100000100000001100111000101110111000100100000011101110010011101110111001001110000011101000111011100100111010000010111010101110011011100010111001001110001011101110111011101110111",
		"01000011011100000111010001100110000001110111011101110111010000000000011100010111000100110110010001110100011101000111011100100111001101110011011101110111001000000111011101110000011100110001000100110110011101110111011001110111011101110111001001110111000100010110011101000000011101110111011101110101011101110011011100010000011100110111011101110111011100100000011100010111011100010100011100110111011100010111011101100111000101110111011001110111011101110110011100110111001001000111011101010111001101010111011101110111",
		"01110111011101110111001101010111011101110111011101110111011100110111000001010111011101110010010001000111011101110111011101110111011101110001011101010000011100000111001001100111011101110111011101010110010101110010001001000111000101110000011000010111011100010011011101110111011101110111011101110000011101110011011100110100011101110111011101100111011100110101011101110110001001110111000100110100001001110111000101110111000101110000010001110111011101110111011101110111011101110110011101100010011100000111011101110011",
		"00110010010101110110011100100011011100010111010001010101011101110111011001110111000001110111011100110111011100110111011000010011010001110010011101000011011101010000011101110001000001110111001001110111001101110000011000110100001001110111011101110111011101000110011101110010001001110111000101110001011101110011000101110101011101110111000000100111011100110111011101110111011101110111011100110111010000000111011101110111000000110100010000100111010001000000011101110111000001110100011100110011010101110111000001110010",
		"01110111010101010111001101110111011101110111000101000111010001110111011101110111001101100111000001010111011101110111010100000100000001110111010101110101011101110111011101010111011101110110010001110111011101000111001101110110011100010100010101110111001001110111011001000010011100000111011101110100010101110000000000100111011001110111011100100101011101100110011101000111011101110111011101110111011101110000011100100001011101110100001101110111011101110001011101110111001100000001011100010011011101110100000000100101",
		"00110111011100010111011101110111011101110101010100010111011001110010011100100101011101000110011101010111010100110110011101010010010001110111011100100111000101110111011101010111011101010001011101010110001100110111010001110111000000100111011100100100011101000111001001110111011100110000010001110111011101110111011101110111011001110011011101110111011101110101000101110010011000000011010100110000011101110111000101110111001001110110011101110100011001110000011100010111011100010111011101110111000001110110011101010101",
		"01110011011101110110011101110111010101110111001001110111011100100111011101110100011100000111011101010010011101000010001101100010001001110110011101110111010101100100010100100110011101110111011101110100011101110001011100000111001001110111011101110111011101110011011101110011001000010111011101100010011101110000011100010111011101010111010101110001011101110000000001100111011101110111011101110011001001110111001100110011010001000000000000000111011101110111000101110101010101110111010001110111011101110111000000110101",
		"01110111011101110111010101110111001001110111000101110111011001000111010001110111011101110011011101110111011101110101011101110000000100010111011101110111011100000000011001110101011101010111010100000010011100000111011001110111010001110001011001110111011100010111011100110111010101110011000001110101001101110101011100000010011101110111010000100111011100010111011101110101011101110111001001110111011101000001011001110111011101100110010001110111011101110011011101110011011001000010011001100111010001010011011101110011",
		"01110111000000100000001101110010000001110000010100000001011100010111010101110001011101110110011001110111011101110111011101110011001100100111010101110111011101010111010001000111011101110001011100110111011101110111011101010000011101110110011100010111001000000111011101100111001001110111011101110010000101100011001001110111000000010000010100110111011100010111000001110111011101110111011001110001011101110011011101010101011101110111011101110111010100110100011100100011000101110000000101110011011100010111011101110111",
		"01010110011101110111011101000010000101110111011101110110001101110011010001110010001100100111011101110111011101110000011100110111011101010111001001110101011101110111011101010111011100110111011101010111011101110001011101110101011100110001011101110111001101110111000101110100011101110010000001110001011101100111011100100111011101110111011101110101001101110000011101110110011101110011010001010111011101110111001100000011001101110111011100010111011101110111011101000111011001110111000001110111011101110111011101010010",
		"01110111011101110111011101110111011101110111001001110101011101110111000100010111011101110100011101110111001001110101011101110111001000110010011101000111001001110111011001110111011101110101011101110111010101110001000001110111011101000111010101110111011101110001011101110111011100110111000101110101011101110111011101110111011001000111011001110111010101110101011101110111011101110111011100100011011101110100001000000111011101010111001100010111011101110111011101110100000001110011011101110000000100110111011101100111",
		"00010111011101010000011100110010011101110111000101010001011100000001011100000100011100100111011101100111000001110111000100100011001001000111011101110111011101110111011101110111011101010111011100110011001101100101011001000110011100010001011101110111011101110010011101000111000101110111011101010110010001110111011101110111011101110111011101110111011001010111011100100110010101010011011101000111011001110010010101110100001001110111011101110111000001110111011101110000011101010111010101000100011101110010011101010010",
		"01010001011100110100010001110111011101110111011101100000000101100001010100000111011100110111011101110101000101110111000001010101011101110110000001110100011101110111011101110111011101010100011101110010011101110110011101110111011101110111010001110111010001110111011101110000011101110111011101100111011001110111011100100111011101010111000000110111011100110010011101110110000001110111010101110000001101110111011101010111010101000111000000110101011101110111011101110001010101110011000001110000011101110111011100000011",
		"01110010011101110100011101110100011101110000011101110101011101110111000100100011011100110111011001110111000001010110000001010111011101110111011101110111011101110111011101110011010101100001000000100111000001110010001101110111001000000111011100000001011101110111001101110111000001110111011100000111011101000111011101000111010001110111011101100111011101110111011101100111011101110100011100110010011100010111000100100111011101110000001001110111001101110111011100010111011101110011011101110111001101110111000001110111",
		"01110100011100000111011101110111010101110111011000110001011101110100011101100111001000100001011101000111011101110111010101110001001101110111010001110100000100000111011101110111011100010111011100010100001001110111000101110111001001110000010000000101011101110110011100000111001001110011011101110111011101110101000000100010011101110110000001110111011101110110011101110011011101010111000101110111011101000111000001000111001001110111010000000111011100010110010001110101011101110010011100000111011101000001011100000111",
		"00110111001001110111000101100111011101110000010101110111001000100111011001010111000101000111010000010011011100110111011100000111011101110111011101110111011100010111011100010111011101110111010001110111001001110111011101110111011000000111011101110010000001110001010000100110011001110111011101000000011101010001011101110100011100010111011101110111011101110111011101110010001101110111011100110111001001110111010001110111011100010110000001100111011101110100011100010000001100000111011101000111011100110111011101110100",
		"01110111010101110000011100100111011101110100011101110111011101110101011101110111011100110111010101110111011101110101011101110111010101110101011101010111011000010000010100110111011101110100011101110111011101110111011100000100011100110110001001000000011101100111011101110111010000100111011101000101001101110111001101110111011101110111011101010111000001110011011100110111011100010111011101110011011101100010011101110111001101110011011001100100010000110110011100010100000101110010011101110110011101110101010001110111",
		"01110111011100010011011101010010000001110100011100010111011101110111000001110111011101110110011101110001011101000111001100000111011000100111011101100111011100100111011100100111011101110110011101110110000001110010010101010111011101110010010001110010001101110000000001110100011101110111011101110000001101100111001100010011010001110111010101110110011001110111010001110100001000010111011101110111011101000110000101100011010001000111010101110111010100110111001101000001010101110111010101110111010101010111011101010111",
		"01110011000001110001011101100111001001100000011101110111011101110111010101110111011100010110011101010111001100100111011001110111011101010111001101110111001101100111001001110000011101110000011101110100010101000100011101110111010000100011011001110111011101110111011101110111011101110100011000010111011101000100011101000100010001110111011001000010000000100111000101110000011101110010000000110111011101000111011101110111011101110111001000010001011101110011011100110111001000010111011100010001011101100110011101110001",
		"01110000010000110110010001110010011101110111001101110111011100110001011101110011011101110011011101110101011101110001011101110111011101110010001001110111011101110111011101110101001001110011001101110111000001110111011101100111011100110111010001110010010000110111011101110000011100110111011101110000000001110111011001110001011101110111010101110111010101110111011100110111000101110111011100000111011101010111010001000110000101110000010101000010011101000111000001110111011101110100011100010111011101110111011101110100",
		"00100010011101110111001000100111011101110111001001010100011101110110000001010101011001110111011101110111000101110101011101110111011100010111010101110010011101110111011101110111011101110111001101110010010101110010011101110111001000110011011101110111011101110001011101110111011101110010011101100111011101110111011101110111011101110100000001110001011100110111011101110000000000010111011101010001011101110110010101000000011101110111011101110000011101110111011001010111010001100111011100110111010001110111011101010111",
		"01000000011101110111000001110010011101110111011101100111011100110111011101110111010101110111011101010100011101010000011101010111011100100111011001110111011101110010001001110110011100000111000001110101011101110111011001000111011101100111011101110001011001110000011100010111011101110111011101110000011101100100010000100111011100100111011101100000011101110100011101110001010101110100011100000011011100110001011101110000011101110111000100110100011100100010000001110001010100110010011101110111011101110001001001110111",
		"01110111001101110111011101110101011101010011011101000111010101110011011101110100011101110111001100100111010100110111000001110111001001110011001101110111011101100111011101110100011101010111001000010101001000110111011101110100011101010111010101110111011101110011010101110111011101100010000101110111011101110111010001110110000101010111001101110001011101110101000101110000011101100111000001110110010001010110001000000111011100000111010100110111000101110111010001110011011101110001011100110111001001110010011101110001",
		"00000111011001110011011101000101011101110000001101110100011101110111011101110000011101100111011101110010011100110100011101110100001001110101000000010111011101110111000001110111001001110010010001110111011000100010011101110100011100000111011100110101000101110111011100100111011101110100011101110111011100000110010000000111011100000010011001110000011101110011011101110110011100100111001001110111000101110110011100100111011101110111000101100111011101110111010001000111011101110111010001110110011101110110011101110111",
		"01000001011100000111011101110111011100010001010101110000010001110111011100100111010101110110001001110111000001000010011101010111011101110111011001110110010001110100011101110101011101110010000001000101001100010111010001000111000100000001011101110111011100000111011101110001011101110111000001110111011100100110000000100111011100100111001000100000011101110000001001110111011101010111011101110101011101000111000001110111011101010110011101100110010000010111011101110111011101110011011100010111001101110001010001110111",
		"01110111011100110111011100110001011100100111001001110111011101110101011101000100011001110111011101110111010101110111000101110111000101110111000101110101010101110101011101110010010101000011001001110111011001110111001001110111010100110011010101110011011100000011011101110100010101110111011101110111001100010011011101010111011101110111011101110111011100000111011101110010011101110111011101010111011101110101011101110010000101110110011101010100011101000111010101110111000000110111011100000101011100010101011101110111",
		"00000111000000010111001101110111011000010110011100000111011100100000011101110111011100010111001001110111010101110100011001110111000001110111010000000111011100010111011101110111001001100100001100100011011101110100011100000111011101110011010100110111000100000011001101110001010101110011011101110001011001110100001001110111010101000111011101110111001101110111001000010111011100110000011001110111011101110111011100010011001101100100011101110111000101000111011000010101011101110000011100000111000001110100000101110010",
		"01100001001100000010001101000111011100110100011101110010001001000000010101110000011100110111011101110111000101100101011100100100011001110111011101110111011100000011011101110111000000010101001001010100011100010001011101010111011101010100011101110101011101110110011101110010011101110111001001110000011101110001010000110111011101110111010101000111011101110111010101110010000101110011000001000111011101110111011001110110001101110111011101110110011101110101000100100100011101110010011101110111010100000111011101110111",
		"00010111001101110111011101110011011100110111011100100111011101110111011101010101011100000101011100000111011101110111001001110111001001110000010001110001011101110101000000000111011101110111011101100010000001000100011101010111001001010111011100010110011100000001011101100111011101000010011101100000011101110101000101110010011101000111011101100110010101110111011101000010010100100111011101110110011101000010011101110111011100000111000000110111000001110011011101110110010100000111000101110100011101000010010101110110",
		"01100111011101110111000001110000000101110101010101110111010100110100011100110111011100110110011100010111011101110010011101110111011101110000001000110111010101110100011101110111001001110111011101010011010001100111011101100111011101110111010001110111011101000110010101010111011100010001011101100111000001110011011101110111011101010000011101100111011101110001011101110111011100010011011100110111011101110111011101000011000101110111011000000001011000110111011101110111011001010100011101000011011101110010001100110100",
		"01110110011101100001011101110001000100010111011101100111011100010111001001110100011100100000011101110111011101110110011001110111011100000111001000010000010101110110011101110101001001110011011101010111011101110111011101110111011001100101011101100001010101110111000101000011000001110101011000010001011101110111011001110011011100100111000000000111010001000111011101010111011101010111000001110111011101110111011101110111011101110111011101110111000001110000011101010111001100010110011101100111010001110111011101110101",
		"01010111011101110001011101010111001001000100011101000111000100010101000001000111010100010001000001100001011101110110011101110111000101100011010100100111011101110010011101110111011101110000011101110111000001110111011101110011011001110111010101100110011101010111011101110100000001110000011101110011011100010111000101110010000101110111000001110111010101100101001001110101011101110110010001000000010101110111011101110111010001110001011101100101010000000010010100110100000101110111011100110111010101110011011000010111",
		"01110111000101110100001001110111000001110111011101110111000001110011011101110101011100100111011101110101010001110111011100110111010101110100011101110111010101110111001001010111011100010001011101000111001101000010000101110111011100100101011101110000011101110001011100000111001000110100011101110111000101000100010000010111011101110000011100100110001001000110011100110111011101110111000001110011011101110011001101110111011101110101001101110011011101110111011101110100011101110111001101110111011101110100000100110101",
		"00000001011100100000011101100001001001110111011101110110011100100111011101110100010001110111011101100111010000000101011100010101011101110001000100110111011101110111011101110001011101010101011101110111011101110111011101000101011101110101011101110111000100010111010000010011011100010111011101110111001001110010001001110111010001000101011101110010000101110111011100010111011101110101011100000111001001010100011101110111011101110011000001110111001101110101001100010111011100100001000100100110011101110101010101100001",
		"01110111011101000001011101110000011101110111011100110111011101110111011101110100010100100000011101110111011100110111010101110100011101000111011001110111011100110110001101110111010100110011010100100111000001010010011001110111010000100111011001110111011100000100001001000101001000100111010100110010011100000000011101110111010001110110011100100111010001100101011100110010011101110111011101110111011101110111001001010111000001110110001000000101010001110111011101110111011100100111011101010111011000000111011100100010",
		"00110100000100010111011101110010001001110010011101110111011101010111011101110111010100110001011101010111011101110011011001100111011100010111011000110100011101010111011101110000011100010110011101110010010100110111010100110111011101110110011101100000000001110111011100100010011101110111011101110001011101010001001001000110011101000011011101110010000101010111000101110111011101110111011100010111011101110111001000110000011100010111011101110000011101110111011101110010010001110001000100010111000001000111011101000111",
		"01100111000100000111011101110111010100000111011000000111011100000100001001110101000001110111000101110101010000110111011101110100011101000111010001100111001001110000011101110100011000100011001001110101011101110000011101010110011000100100001001010111011100000110010100000111010101000111011101110000011100000001000101110000011000110111011101110110000101110101011001100111011101110111010001110111011000110001000001110111011100000111000101110111011101100111011001110011011101110000011100100000011101100111010001110111",
		"01010001011101110111011001000111011101110110000000100111011000010111011101110100011101100100011101100111000100110111011100100111011100100101011101100111001100100111011101100100011101010111011101110111011100000001011100100111011101110111000000110101001101010111000101110011000100110111011101110111011100010011011101110011011101110111011100100001000000100010011101110110011101110001010001000010011101110100001000000111011100100000011101110111011101110111010001110111011101110011010101110001011100010111011101000001",
		"01110111010001000011010101110111011100110100011001110111011101110111010100110110011101110000011101110111000101110111011101110111010101110100011101110111010101110111000101110010000101110111011100000000000001110011011101110110011001110011010101110111011101000111011101110111011100100100011101110111010101110111001001000111001101110101010101100110010101100000000101110000011101110111011100000111011100000111011100010111010000000011001000010000011001110101011101110111011101110111011101110100010101110111000101110001",
		"01000101011101110111011100100100011000010100011101110111001101110010011100100111011100000111010000100111001000100111011101110111000000010111010101110111011101110111000001110111011100000010011101110111011001110111011100000111000001110011011101110111000101000111011101110110011101110111011001110111011100000111011101110100011000010010001000110100011101110111011100110000001001000011011100100111011101110111011101010110011101110111011101110111011001110111011101110111011001110100011001010011001001110111001100110110",
		"01110111011100110010001100110111011101110100011101010111011001110010011101100111010001110101011101100111011100010000011101110111010001110111011101110111000001110011011101000111011101110111011101110111011101110111001000100000000001010101011000000000000000100110010000100110011101010011011101110010011100000111011101110011011001110000011100000110000101110001011101110100010101110011011001110111001101110111000101110100011101010111001001110001011100000101011101110111000101110000001100100100011101110111010100110001",
		"00100010010100000001010100110111011101110111011101110001011101110000011100000111011101110011011101110011011101110111001000110100011101110001011101110111001001110111011101110111001101110001011101110100011101110111001101110011011101110111011101110101010000010111010001110111011101100111011101100011011101110111011101110001010101110101011101110111011101110111011100100010010101110110011101110010011101110010011101110111011101110111011101110111000100100111011101100011011101100001011100100010000101110101011001110111",
		"00000111000101110011000001110111010101110001001101110100001101110111010001100111010000000111011101110110011100110111011100000110010001110111001001110001000001110010000101110111000001000110001101110111011101110100010001110011011101110010011100010101000001100010011001110111000100110100000101010111000101110111011101110111001101010111011001110111011101110000010101110111001100110101000000000001010001110111001101010111010001110101010001110100011101110111011101110000011101110111000101100111011100000111011101110111",
		"01110001011101110110011101110111011101110001011100110111011101110111011101110111000000010111011100100101010001010111011101110111010000110100011101010111001101110111011100010111001001110000011001100100011101110111011101110111000001110010011100110101011101110110000101110010011101100111000001100011001101110010011101100111010001110111011101110111011101100111001001110111011100110111011101010111011101110010010001110101011100000111010000110100011101110111011100100001011101110111011101010111011101010010011101110111",
		"01110001011101110000011101000111011000010111011101110111011101110111011101010111011101110000011101010101011101000011011100010111011100000111011101110111000101000101011101110001011101110100011101100010010000010100011100100111010101110111011101110111011100110111010101110111000101110100001101110110011101110111001100000111011001110111011101110010011100010111011100010111011101100100000101010111011101110111011101110011011101110111011100100101010101110111011100010111011101100111011100000111000100000110011101110111",
		"01110111011101110100011100010111011101110111010001110111000001100110011101000001011101110111011101110111010100100111011101110111011101110111011101110111011101110111001001110111011100110111011101110000001001110111010000010111011101110000011101110011010101000001010101110101000100100111011001110111000100000101000101110000011101110111010100110111010000100111011100110010011101110010010001110101000101110111011101110111011101110111011100000101011101110111011001010111011100100111011100000001011100000111011100000110",
		"00010111001100100111011001110111011101110000011101110010011101110111011101100101011101110111011101110111011001110111011101000010000001110111011101100100000000010010011101100011001101110010011101110111011101110111001000010111011100100010000001110100011101110010011101110111011101010111011101110010011100100010011101100000011101110001001001110010000001110111000101000000011101110100011100100101011101110001011101110011010100000111011101010000011101110111010100100111001101110111011100110111011101100001001001010111",
		"01110010011101110111011101100111011100000111011101110001010001100011011101110001011100110101011101110010011001110111011100100111000101110111011101000111011101110000011101110111000100110111010001010111011101110110011101110111011101110111011101010011011101110010011101110100011101110001011101010011011101100111011100110101011101010100011100110100011101110010011101110110011101110111011101110111011101110111011101110110011100000111001101110100011100100101010100110111001101110111011100110111011000100111011101110010",
		"01110010011101010111010001000111011101010111001001010111011101110111001001000101001001110111011101110111011001110000011101110111011101110111011101110110001001110111011101010111011100000001000000010111011101110111010000110111011101110111011000100100011101000111010100110111010100100001011101110111000101110101011101110111011101100111010101110111011101110111001100010001011100000111000101110101010101110101011101110111010100000000011101110001011001110111011100100110010001110010011101110100001100000000011101110010",
		"01110001011101110010011000010111011101110110001001110110011101110011011100100111001001110111011100000111011101110111011101110111001000110110011101110110011101110111000101100110011101110111011101110111011101110111000000100111011001110100010001110111000001110010011101110100000001110111011101110111000001110111011100110100011001110000000000000111001001110111011101110111011101110000011101110111011001010111011101110010011100000111010001110111011101110101001101110111011101100100010101110000010101110000011101110000",
		"01100111011101100010011101110111000001110111011101100011000001110111010101110010011101100111011101110010010001110100010100100001011100100000011101100000011101000111010101110010011101110100000101110000011100010111011101110100011101010111011101110101011100110111011101110010000001000111011101110001011101100111011100010111010001110111010000010111010001110111000001110111010001110110011101110111001001110000000101110111011101110110010001110111011101110000010001110111011101110111011101110001010101110010011101010101",
		"01110110011101110110011001110000001001110001001101110111011101010111010000100111011101110111011100010111011101100111000001110111000001100111000001100111011100100111010101110111000101000111011101010111011101110010011000010111011101000111011101100011011100100010000101100111011101110111011101110011011101110111001101110001011100110111011101100111011101110111001001110110011100100111011001110111011100000010001001100010011101110111001001110111010101110111011101110111011101010001001100110111000001110010011101110111",
		"01110111011101110101011100000100011101110111011101110111011100000111010101110101001100010111011101110101011101110101011101110111011101110111011100000111011101000111011101110010001000100111011100000010011001110111011101110111011101110101011100010110011101110100000001110101010101110111011101110111011100010111001000110010011101000111011000100011010101110111011100000001000101110111010101110111011101110111001001110110010001110010011101000001011101110110011101010111011101110001011000000101010101110111011100010111",
		"01110111011101010110011101110111000001110111011101110111001001110111011101110111000000000111011100010111011100110111011101110000011101010111011100000111010001110111011101110111010001110001011100110111011100010111011101010111011101110001011101100101000100010111001101110111011101110111011101010111010000010101011101010111011101110111011001110111000100000000000101110111011001110111011101110111011101110111011000110111011100100111011101110111000101110111011001110010011101110010011000010111011000100111011100000111",
		"01000011011100100111011101110111000001010110001001000111010101110111011101110001001101110000000101100111011101000001011100110111010000100010011101110111010001110111010001000111011101110001011100010100001001110111001000100011011101010111000101110101011101110111011101100111000101110100011100000111000000110111011100000101011100100000011101110111000000000101000001110011001001110001011101110111001000110010000101110111011101110111011100100011011101100111011100010111010101110111010001110111011101000011011101110111",
		"00100100010100010001011100010010011100000110001101110000000101110111011100010110001001110101001001110111000001110111011101110101011100100001010001110010010101000111011101110000011100110111011101110001011101110111010000000111010101110111010101110111011101110000000001110111010101110011011100100111010101110100010101110111011101110001011101110111011101110001011100010101011101110111011101110111011101110011011001110000001000110111011100100111010001110001001101000111000101010111011001110111000101110100010101110111",
		"01110001010101110101011001110111011101100001000001110111001101110011000000010111011101110001011101110111011001110111010101110111011101110011011001110000011101110111001100110111011100100111011100110111011001110111001001110100011100100111011101110010011101110111000001010111011101110101011100000101001001000111011100010101011101110011010000100011011101110000011101110111011101000010011101110011000001110111011101110100011101110000011101110111011101010111011101110101011101110111011100110111011100110100011100010111",
		"00100111011100100111011100100111001100010111011000100111000000000111011101100111011101110111011101110111011101110101011101110111010000100111011100010100001101100110011101110111011100110111011101110101011101110111010001110111011101110010011101110011000101110111011100110010010101110001000001100010010001110111011101010111001001110111011101000111011101010101011100100111000001010111000001110111000000110111011100100100011100100111011101100111011101110010011101110110011100010101011101000111001001110111011101000111",
		"01110000000101100101011101110011011101110111011101110111000101110110010100010100010000110000001100100000000001110011010101110111011101100111011100110101011100000111011101110111000101100011011101010111001101110100011100100010000001110111001001000111011101110111011101110111001000110111011101100011011101110101000001110110011101110111011101010111011101110111011000010111011101110111010101010101011100010111011101110110011100110010011101100111011101100111000101110110011101110110000001110101011100010001011101100010",
		"01110111011101100111011100000100011101110111001001110111011000100010011101010111011101110111001001110101011000100010000101110111011101110100011101110111011101000111000001010101011101110110011101110100011101110111011101110001010100100100011100110100011001110111010001110111011100000110011101110111010101110111011101110111011101110001011101110111001000110100011101000111001101110111000101110111011101110111011001110111011101110101011101110111011100000101011101110100001000000000010101110111011101110111011101110111",
		"01110010011101110111011100110111011001110011011101110111011101110001011101000010000001100111011101110001010101110000010101010111001101000111011101110111000001100111011101110100011101110010011100010111001101110111001000110011011100000101011101110111011001110111011101110111011101110111011001110010011001110011011001110111011101110110011101110111011101110011011101110111000001110111011001100111011100100111011101000100000101110111011101110111011100110000010100000111010001110111011101110110011101000001011101110000",
		"01110111011101110011001100110111001101110111011101110111000001110110011101010111011101110111000100110000011101110111011101110111011101110010011101110001000100100011001001110110001000100111000001010111000101110111011101110111010000110111010000010011011100000101000101110110011000100000000101110010011101110100011101110111011001000110011101010111011101110101011100000011001100010111011100000111011100110001010101110100011101100111011101000100010101110111011000110101011100100111000101110000011101110111001101100001",
		"00110101011101100111011101110111010101010111001101110101011101110111001101110111011101110110011100110101011101110111011101000111001001110100011101110110011101110111011100000111001101000010010101110001011100100111000001110110011101110111011101110111001000010111011101110111011101110000011101110111011101110111011101100111011100010111001101110111011100000111001001110111011101110111011100010111011001100000011101110100010001110110011101110111011100110111011101110010011100110100000101110111011101110110010101110000",
		"01110010011101110001010001110011011101110011011101110111011101010111011101100111010100000111011101000111001000000111011101010011011100110001001101110001000001110111011101110110001001010011011101110111011101110000011101010111011100010111011101000111011100110111011101110111011101010011011101110111011100110111011101000111010001110111011101110111011101110111011100110111011101110001010000110111011100100000001101110111011101100011011100110000000001110100011100010111011100010111011101110111000001110111010001110111",
		"00010111011100110010011101010101011101010110000001110111011000000111000000010111011101110111011101110111011101000001011101010111011101000000011101110111011100100001011101110000011101000111010001010000001101110111011100100111011101110111011101110111011100110111001001110000011101110110011100010111000001110111011101010101000001110111010101110111011101110111010101110111011001110001011000100101011101110001011101110111010101010111011101100111010000100111011101100111010001110111011101110101011101000111000101000001",
		"01100100000101110101011101110011001101110111011101110001011101110110000001110111000100100111011001110100011001110100011101000001011101110111011101110111010000110111000001010111011101110011011101110110010001110001011101000111010101110111010001110111011100000111011101110111011101110111001101110111011101110110011101000111011101110111010101000110011100100001011101100111011100110111001001110111001001110011000101000001011101110111000001010100000001110101001100100111011101010111011101110111011101110111011101110110",
		"01110001011101010111011101110101011101110111010101110100011101110111011001110111011001110111011100010100000101110001011101000111010001110101011101010100011101010111001001110111011100110111011101110111011100010111011101110111001101010111011100000111011101110010010100000111011101110110011001110001001001000111011101110101011100110111011101110110010100010000010000100001011101110000011101110111011000000111010101110111001101110110011101000111011100110110010001100110000000000111011100110111011101010101011101010101",
		"01100111011100000000011101110000001000010111010101110001011101110111001001110101011101110100011101000110011101110111011100000111010100110001001100100110010001110101011101110111011101010111011100010111011101000111010101110111011101110110000000000111011101110111010001110011001001110110000100010111011101110111000000010111011100100000001101110001011100010000011001110100011001110111010100100100000101110101000101110111011100010111000001100001011101110011010100110111011101110111000001110111011100100111011101110001",
		"01110111011001110011011101110111001001110110000101110110011101000111011101110111011101000111011101110111011101110000011001110111000001010111011100000111011101110010011100100111011100000111010001110111011101100111011000010111011100010111001101110000011101110011011001110111011100100111010101110111011101110011011001000111011001010111011101110111011101110001011101100111000101100011000000000001011100000000000000110110001100010111011101110000011001110111011101110010011101110111010001110111010001110100000000100000",
		"01100111000101110111011100000011010100110111011100000001011101110111011101110111000001110111010000100111000001110101011101110111001001110011011000000111011100010111000101110111011001110010011101110001011001100111000101110100011101100111011101110111011101110111011101110110011100000101011101110010011100010111001101110111011101110110011101110011011101110100011101110111011101100111010001110111011101110111011101110111011101010111001001110001010100000101011101110011011101110011011100100111011101110111000001100000",
		"01110111011101000001011001110010011101000001011100000011001000010111001001110111011100110000011101010111001101000000011101100111000101100111011001100111011101100111011101110110000101110111011101100101011101110000011101110111010101110110011101110111001101110111001101100001011101110111001101110111010001110111011101110111011100110111011100000010001001110000001001110111011100010111010101110111011001110111011101010111000101110111011101110000011100110111011101110001011101110001011100100110011100000111011001100111",
		"00110111011101000111011001110101010001110111000001110101010101010101011101110111010001110100011101110111011101110101011100000110001101110111010100110111010000100100011100100000011101010111000101110011011101110111011101000111011100010111001101110111011001010111010101010111010001110110011101110100011100000101011101110010011101110111011001110111011100000101011100110111001001110110011101110111011100110010000101110001010100100001011101110111001000100111011101000111011101000011001001110111001001110111011101110111",
		"00110111011100110111011101110111011101010001011101000111011101110111011101110100011101100111011100110111010101110001011101110100010000100111000000000111000000100111001000000111011101100111011100110110011101110101001000000111011100000111011101110010001101110111011100110010011101110111011100110111011101110111011101110111011100010111011100000011001001110010010001110111000001110001011101110111011100100111011101110100001101110101011101100101011101000111000001110111001101110111011101000100000101010111011101110001",
		"00100101011101110111011101110110011101110111001001110000010101110111011100000111011100000000011101110111011101110111011101110111000100100011011101110100011101110110000001110011000001100000011101110111010101110000011101110100011101110111011100110010011101100111011101110111000101010001011101110100000001000111011101110111000000110111000100100000010101100111011101010111010101110100011000010111011101110111001000100111010101000111011101110111000101110111011101000011011100100111010101000010011101110111010101110100",
		"01110011000101110111011101110111011100100111000101110000011101100111010101000111010101110111010000110111010101110101011101110111001101110111011100100101011101110111011100000011011101110111001001110111011101110111001101110111010001110100011101110111011101110000010000000110011100010111011000100111011001110111011001100111011101000000001001000100011100010111011101100111011100110011011100100110011100100110001101110111011101110111011101100111010001110100011001110100000101110111011100110111011101110011010000010111",
		"00100111011001110100001001110111011100010111000101110111011101110111011101110101011100110100010000110001011101110001011100000111001000100111011100000111011101100111011100110100011001000111001001110011010000100111001101110011011001110111011101010111011101110010011101110100011001010111011100010111000101110000011101110111011101000110011100000111011101010111011001110111011101110111011101110111011101110111010101100111011001110111001001110000000101110111011101110111011100000000011100010111000100010111001001110111",
		"00000111011101110001011101110111011001100111010100110000001101110111001101110101000001110111000101000111010000100011010001110001001001110111010001110111011100010010011101100111011101010110011100010101011100100111001001110111011100000110011100000011011101110111010101110110011101110100011101100010011101110100011101010111001101110110011101000111011101110101010101110011001001100110010001110110010001110111001101110111011101110001001001010111011101110111011101110000000001000001000001110111010000010111011101000110",
		"01110111000001110111011101010111001101110010011101110100001001010111011101110111011101110111011101110111001101110111010001100010011101100000011101110000011101110111011100000111000100010000011001110111011100110010010001110010010101100000011100010010011100100110000001110111000101000111001101110101011100110111011101110111000001110111000001110111000101110001011100100111010100000010011101110111011101110110011101110000011101110011011101110111000101110111011001000010011101110111011101100101010001110000011101110111",
		"01100000011101010111011001110111011100110010011101110111011101110111000101110111011101100111011101110100011001010111010100110111001001110010011101110110011100010111011101110111011001110100001001010111011101110111011100100011011101110001001101110111001101110110011101100111011001110111010101110110011101010011011100010110011101110111001101110111011101110000010101110111011101110111011101010111011001110111010000110011010101110110011100000111011101110010000001110000011001010111011101000000011101110110011101110111",
		"00010101001001110101000001000111011101010111000001110111011100110111011100100011011101110111011101110001011101110111011101110101010101110011011101110111011101110111011101000011011100010111011101110001000001110011011100000010010001110111001001110101000100100111011101110111000101100101011000110111010100010100011100000111010000110111010101100001011101110111001001110111011101000111011101110111000001110111011101100111011101110010000001110110011100100100011101110001000101110100011101110010011101110111000101000111",
		"01010111011101100111001001110001011100010111000101110111001101110100010101110010011100110000000100100111000101110100011101110011011101110111010100010100000101000111011101110110001101000001011101110011011100110100011100100011011101000111011101110010011101110111011100000000001101100111011101000011011000000111011101110111010001110111011100000111001101110101011101110100011101110001011101010111001001110010010001110001011101110001010001110111011101110000010100100111011100010011011101010111010100000111011101110001",
		"00100111011101110111011101110111011101110111011101000001011101110011000101110111000101110111011101110111011001110011010100010111011100100011001000100111011100010111011101100100001101110111011101110111011101110110011101010111010101110111011100010111011100100111011101010111011100010111001001110101001101110111001101010111000101110111011101100111001000010010011101110110011101100111011101110111000101110111011101110111011001110000000101110111011101110001001100100001011101110011011101110101011101100111011101100001",
		"01010111000001110111011100010000000100100101000101000000000101110111001001110000010000110011011101000001011101000110011101110111011101110111011100110111011101000111011101100111000001110000001000000011011101110111001000000101011101110110001100110111011101110111011101000111011100110111011101110111000001000011000001110000010101110111000101110011011101110011011101000010011000100110000001110111011001110000010001110101010001110110011101100111011100000111000001100111010100100111011101010111001100100011011101110111",
		"01110000011101000101011101010010011101110111011101000010011100100100000100110111011101110100011101010000001101110111010101110111011100110100000001010001011101110101011101110111011101110000011101110101011101110111000101110110011101110111000001000100010001110111011101110001011100000111011101110001011000100001011101100011011100100100011101110110011101110111000101110111000101100101000001110001011101110111010001110000000001110011001100100111011101110110000001110101011101100101001001110111011101110110011001100110",
		"01110001000101110001001000010001011101110001011101110011001101000111011000100100001101110001010001110000000100100111001000110010011001000111010001110101011101110111011001100111010001100101011101110111011101110100011101110111010001110001000101110111011001010000011100010000011100110111001001110100011101110111011101110111001101100111011101110111011101100011000000110110011100100000011100010111011101110011011101110111010001110100011101110011011101100001010001110111001101110100000001110111011000110111011101110111",
		"01110111000100000101011101100111011100000111011100110111011101110100011101110010011101100111011100100111010001110001001101000111011101010111011101110110010001010111011101110101011101110111000001110111001101110000011101110111011101110111011000100111000001110111011001110110011101000111011100110111011101110111010101110111001001110111011100110101010001110010010001110111011101110001011101010101011100110110001001110111011101010010000101100110010101100010011101100111011101010111011101110011000101010111011101110111",
		"01000000001001110111011101110101011101000111011001110111011100110000011101110010011000010111011101100100010101110111011101110111011100000010011100000010001100000111000001000111011101110010011101110111011101110111011101010111011000110110011100010110011101110111011101110111011100010000011101110111011101000111011101110111001001110001011101110011011101000111001001110111001100100010011100110110000001100100011101110100011000010100011101110111011100000111010000000010011101110010011101110111011000100000011101110111",
		"01100111011101010111011101110111011101110111011101110110010000110000010001000111011001110111011100010010011101110111011100110000000001010111011100000001011101110111011100000101011101110111011101110111010101000010011101110111000101110111000101010111011101100111010001110111011101110001011101110111011101110011011001110001011100100111000101100011010101010111011000000111001001000100011001110101011101110111011001110111011101110000010101110111011101000101011101110111011101110111000001100000011101110010011001110111",
		"00010010011101110100011101110111001100100010011101110111011001110111011100110001011101110111001100100001011101110111011101110111000001110111011101110100001001110001011101110011011100100111011100110111011101110111011101110111011101110111000001110111000101110111011101110111011101110111011101000000011001110111011101100001011101000111011100000010011100000101011101110100011101110011000001110111001001110111011100010111000101100111011101000100011101110100010101110111011101100111011101110111010101110111011101100100",
		"01110011001000110010011101000111011101110001001001110001011101010111011101010011000101110111011100110100011100010100001001110111011101100011001000000111001001000111011101100011010101110111011100100001011101100010010101010111011101110011011101110001011100110101011101110111000001010101011101110000000001110100011100110101011101110111011100010001011101110111011001110111011101110100011100110001001001110111001000100111011101100111010100110111010101110111001101010001001000100111011101110011001101110111001001110111",
		"01110101010100110111011101110010011100000111010000010000001101110100011101110111001101110000001101110111001100110100001100010011011101110111011101110010011100000111011101110011011000000111011101110110011101110111010001010100000101110101010001110111011101110001011101110111011101100111011101110111011100100001011101110111011001110111011101110011011100110111000001000010001001110111011100010111001001110110011101110001010101110000011100010000000101110101001101110101011101000001011101110001011101110100000001000111",
		"01110100010000000111011101110000011001110111001001110111011100000111011101110111001101000000011101110111011101110000011101110001010100100111010001110111010001010111011101110111011101110101000000110111001101110111011101100111011000010011011100010110011101110111001001110010011100100000011101110100000001110111010000010111011101110111000001110001011101110111001100100001011001010011010001110101000101010111011101110111001001110111011101010111011101110100011100100111010101110111011101110100011101000111011101110111",
		"01000111011101110111000100010111010101100010010101100111000101110000011101110010001101110111010101110100000001110110011101110110011101110011011000100101011101110001011101110111000001110111011100110100001001110010011101110111001001010111000100000111011100110011010001110111000001110111011101110111011001110111011101110111011100100001011101110111000001110001010101110001010000100111011100000101011101110001001001110111011001110111011101110100010001110111011101110111011001010011000100000111011100000111011100100111",
		"00100111000001110010001100100111011101100001010100000111011101010111011000010111010001110000011101110000011101110100000101010010011001110111011101110000000101110100011000010111001000010101011101110111001101110111011101110000011101110111010001110111001101110101000101110111011101110101001001100111011100110011011101110111001100100111011001110101011100100111011100000111011101010111011100000111011100100111010001110010011101110110000101110111011101000111001000010111011100100111011101110111011100100100011100110111",
		"01110011011000100111011100110111011100110111011100100001011101110000001100010010011100100111011101110111011101110111011001110111001101110111010100110101011101110001011100110101011101110100011100000001000001110100011101110111011100010000011101110111001001110100011101010111010000100111000001110110000100110111011101110110011101110111011001110110011001000110011101110000011101110111001000000100011101110011001101110000011100110111011101110111000100100111011101100100011101110111010000010101010100100001011100010011",
		"00000111011101110111010101110110010001010101011101110111000101110101001001110010011101110111011100110111011101110000011001110001011001110010001100010101011100110110010001110111011101110101011101110001011100110111000101110111011101110011011101110111011000000111011101010111001001110111001100010111010101010111011101110001011100000000000001000111011101110000000001100100010100110111011100010100000101110101010001110111011100110101011001110100001001110000000101110111011001110000011101110111010100110111011100110111",
		"01110101010001110111011101110111011101100111011100110101000001000111011100000111000101010111011101110100011101110111001000010111011101110001000100110110011101100111010101110000011101110110011000100111011101110111011001110111000001110101011100000000011101110010000101110111011100100111011101110111011101110111011101110111011101100001011100100111011101110111001101100101011101110111011101110111011101110111010001110111001101110111001101010001011101110111000001110111011101110010000101110011011101100010011101110010",
		"01100111000001110001001101110101001101100110010001110111011101110011010001110111001000000110011100000001010101010010011100110111001101110001010101110111011100100111001101110111000101110110011100010101011101110111011101110110011101010111001100000111011101100001011101010011011101000111011001110000011101110110011101010111011101110001010001110011001101110110010000000100011101110010011100010101011100000100011101110111011101110111010001010111011100000111000101000111011001100100000001110000011000000010011101000011",
		"01110011000101110111010001110111010001110111001100100010001001110101001101110010011100010000011101100111010001010110000100010100011101000111001001110011011101110111010001110111010000110010011001110101011101110111011100110001010001110110001101010000011101100111011100010111000101010100011101110001011101110011011101110010011101110111011101110111011101000000010001010010011101010111000100010111011101110111011100010011011101110111011101110001000101110010011100010001001101100001011101110010011101110011011100010100",
		"01010101011101110111001001100111011101100111011101110111011001010111010101110101010000000111010001110111011100000111011101110000011100000110010101110001011001110111000001110001011100100111011101110111011100110111011100000011011101110100001101110101011101110111011101000010011101110101011101100101010001110000011101110111000000100101010101100100011101110111011101100110011100100010010001110000011101000111011101110111011001110010011100100111011101110111001000000101011101110100011101110110011101110101000001110111",
		"01110111001001110100011100000111011101110111011101110111011001010111011101110000011101000010011101110111001000000111011100000111011101100111011101110000011100110111000100100111011101110100000000000010011101100111011101100110010101010011011101110111011100000000011100000000011101110111010101110111011100110101011101100111000101110010010001110111011101110100010100100111000101110111001101110010011101110100011001110010001001110110011101110111001101110010001101110111010001110111011101110111011101110111010100010111",
		"01000111000100100100001101110010000101110111001000000111011100000010001101110010011101110111011101110011001100110111000001110011011101010111011001110111010001110011000101110001011101110010011000100111011100000111011101110110011101110001011101110111001101110111011101110111011101110111000000010111011101110100000001110111011101100111011100000101011100000011001101000111011001110001001101100111000100010111000101110011001100100100000101110000011101000111010001110000011001110111011101110101000001100111001101110111",
		"01100000011101110111011101110011011100100111011001110111011101100110011100000000001100010111011101100111011101100001011101110111001001110111000101110111011001100001000101110111010000010111011101110111011001010111011101110000010101110011000001100111010001010111001001000110010101110111010101110111011101010111011101100111010001000111011101110111011101110111011101010111010001110111001101110000011101110111000101110111011101110111011000100111000000100111001100000100001101110111010100100111000000110101000001110111",
		"01000111011101110100011100000111011000100111000101000111011100100111011101100111011101110010001001110111011101100111011101000100001001000001011101110111010101110011011101000010011101110100010001110111011101110010011001110111011100110111010001000111011101110111001101110111011101110111000001110011011101110001000101110111011101110011011100010111000001110111011101100111001001000111001001010111001001010111011100010110011001110111000101110100010101110100011001110111011101110101001001110111011100100101011101110111",
		"01110001011101110100011101110111001000100000011101110110010101110011011100000111011101100011011100010100000001000111011100010011011000110111011101110010010100100111010001110111011101110100001101110110011101100111011100100001011101110010011101000010011101110011011101110101011001110111010001110101011101110100011101110111011001010111011000000111010100010111011101100111011101110111011101110111001100010111011101110101011100100111011101110111001101000111000101110111010001110111001001110111011100010111011101000111",
		"00110111011101110111011101100111000101110101010001110000001101110100011101110001011100110111010001110010011100000011000101110001001001100001001001110110010101110111001000010111010101110111011100000111011101110111011101110010011101110111011101110100011100010110011101000111011101110111010101110111001000100111011100110010010100100111000101110000011101000111011101110111011101110111011101110100011101110110011101000111011101110111011101110010010100000111011101000001010001100110000101110111011101110111011101100000",
		"01110111011001110000011101010111001001110111011101110111010001110000011100000101010101110111011101110000000101010111011101110111011101110111011101110011011101110001001100010010000001000111011101110110011101110111001101110011011101110101011000100110010001100111011101110011000001110111011101110100011100010111011101110000011101110100011101110111010001110011011001000000001001110010011100100111011101110111011101110011011100000101000101110111001100000111001101010111011101110111011100110111000101000111010001110010",
		"01000111011101110111011101110111011101110110011101110111011101110111000001110111011101110111011101110100001001110100011001110010011001110010011001110110011001010111011100110111011101110100011101000111000001110000000001010111001101110111011101110010011100110111000101110111011101100011011001110111011101100111011101110010011001100101000100110000011101110111011101110111011100100111011101010111010101110111001100000001011101100000011101110111010000110111011101110100000001110111000000010111011101110001010101110010",
		"00110010011100110100011101110010011100100111011101110110011101110111000101100110001100010111011101110111011101110110001001110011010101010001001101010111011101110111011101110111010100000111011101110111011001110111011101010110001101110101011101010111010001010100011101100011010001110100011001110100001101110111010101100111001001000111011101110111011100110111010101010111011101110001011100110101001101110111001001110101000001010111011100000111010000100100011101010111010101000011011100100111010101000111011101100100",
		"00110111001001110101011101110011001100100111011101000111010001110111010001110110011101110111011000100111001101110011010001110111011101100001010100100111010101110001011101110010010101110111010100100111011101110100011101110111011101110111011100110111000101100111011101110111010101110001001000000111000100000111011101000101001100000111011101000000001101110001011101110101011101110010011101110111011100110110010001110011001101110010011101110111011001100100010101110010001001110100000101110000011101110111011001000000",
		"01110111010101110110010000010111011101110011000101110110001000110111001100110000010000110100001101110111011100110111011101010111011101110001011100110001011001010111011101110111001001110111001101000010001001110111011101010100011101110111001100110000010001110110001001110111000101110111000001110010001101110111011101110111011101110000000101110111010001110111011101110111011101110011001000100100011101010111011101100010011101110100011101010111011101110111011101110111011101110111001100100001011000100010011100100111",
		"01100011010001110111011101110111011001110111001001110111011101110111010100100001011101110111011101000111011001110111011101110101011101110111010100010101011100100111000101110110011000110000011101010111011101110011011101110111001000000101010101110001011101110001011101110110000001100111011101010111010001110111011101110001011100000111011101110100011001110111011001110000000101110000000001110111011101110110011101110111001101110111000001110011000001110111011001110111011101100111011101110111011100010111011101110111",
		"01100111011101000111011101000111010100100111010100010111011100110111000001110000011001100111010000110100011101110100001101110111011100100101010001000111011100100111011101110111011100110111011101110100011101100111011101110111011101010111001001110111011001110111011000000111000101110010011100100111011100100111000100000111011100100111011101110000000001110011010101110111011101000000011000000101011101000111001101110111001001110111011101110111010100110111010101110110010000000110011101110111010101010010011100000110",
		"01100111011101110001011101110110010001110111010001110111011101100101011101110111001001110110000001110101011101110111010101110111011101110001011101110100010101110010010101010110011100010110000001100111011101110111011101000111011100100111010101110111010101110111011100100011011100000111011101110111011101010001011101010111011101110111011001110101011101110000011101010111010101110001010101110001011101110101010001110111011101110111001101110111001001100111011101110100011101010011010101110001001100010010011101110111",
		"00110111011101110101011101100111011100100100000001110101011101010000011101110101001101110111000101110111010000110011011101110111010101110010011101110111011101110111010101100111011101110111011101110111010101110101000001110001011101110001011101110111001100010110011100000111011101110111011101110000011101110000011100100111011001100010011100010110011101010011011101110111011101110111000100110111001101110101011101100011011101110100011101000111010101100111001001110111010100000111000101110111001101110111011001110000",
		"01110111010000100111011101100111011101110100011101010111001101110110011101110111011001110111011001110101000001110100011101110011011101110100000001110001010001110111011101110110011101110111011100100110011101110111011100110111010101110111010001110111001001110000011101110111000101000111010001000111011101000110011100010001011101110111001101000011011001010011011101110110011101110111010001010111011100110111011101110111001001110111011100110111010101110101011101100100011101110111011101100101011100100111001101100111",
		"01100011011101100111011001110101001001110111011001110010000101010110000101110111000101110111011000010001011100100000001001110100011101010111011100100101011101110111011100000111000001110010011101100111011101110100001000000011001000110110011100110111011101110111011101110000011101100111000101010010000001110111011101000111000001110111010001110111011100000111011101110111011100100111011101110111011001110001011100110001011001100111011101110111010101110111011101110100000101110101001101110111011100110101011101110011",
		"01110010001000000111011101100111000101000110011101110111011101110100011100000100000001110011000001110000011100010111011100010100011101110111000001110100011100110111000100100110011101100000011101110111010100010110011101010111000101110111010101010111011101110000011101110000011101000111011101110111011100100111001101110111001101110111000001100111010100000111010000010111011101100000010001110111001001100100011101110111011101110111011101000111011101110110001000000011011001100111010100100000000000110111011001110111",
		"01100110011101110000001101010111011100010000001001110111011101110111001100110100011100110011011001110111010001110011011101100111011100110110011101010011000101110111011100100111011101110100011101000000011101110001011101110100001001110111011101110110011001100101011100010001011101110111011101110111010001110011011101110111011101110111000001110111011100110100001001110100011101110110011100100010010101110111011001110111000101100011000100000111001101110111011101010101000001110111011101110000000100000100000000100010",
		"01110110011101110011011101110100011001010100011100100101011101110010001101110101011100000111011101110011011100100111011101110111010001110010011101110110010001110101010100000010000000000100000001110111011101110010000000010111011101000101010100000111011101110001011101110111011101010111011101110110000001100111010001110101011001100011011101100010011101110011011001110110011100000100011101010110011101010110010101110111010001100111011101110010011001110111000001110111011100100111000000000001011001110000011101110101",
		"01110111011001110110011101110111011101110110000001110001001001110111011101110111000100010001011101110111000101000111010000110101011100010010010101010000011001110111011101110010011100100000011101010110010001010010001100100111011100110010001000110000011101110110001101110110011101110111000001110111010001110010010000010111011101100111001000000101011101110111011101110011011100010111011101110100010001110111001001100110011101110111001001110111011100000111000101110000011101000111011101000011011000110111011101100111",
		"01110111011001110111010000010110011101110001010101110111011101110111001001010111000101110111011101110110011101110011001101100111001101110111011101010111011101110111011101110111011100100111000001110111011101110001010101110111011101110000000101100000011101010111010001000111011101110111010101110111011101110111000101000100010001110010011101010111011100100111011101110111011100110110011100100111011101110111011101110110011101110111011100110110001100110111000101110101011101110110011100100011010001110111011101110111",
		"01000001011101110111011100010111001101110111010100100111011101100111011101110111011101110111011101110111011101010111010000010101011000010001011101110111011100000000010001110101001001110111000101110111010100100111011001110111011100000111011001110011011101010001011101110111011101110111011101110000000101110111001000100110011000000110011101110111011100100100011101110111010001010111011101110111011100000111011101110111011101100100011101110111001101000111011101110111011100000001011101010011011100000111001001110011",
		"01110110001100110111011001010111011101110100011101110011011101110110011101100100011101110111000001110111011100110111010001110000000000110111011101100010010001000111011101110111001001110010010100110111011101110111011100010111010100000111000001110111011100010111010101100100011101110111001100110001000001110111010001110111000001110111011101110100000001110111011001010001010001110100011101110111011101010010011100110011011101110111011101110111011101110111000000000111010001110111000001110010011101000111001001110111",
		"01110111011101110111001101110111011101010100011101100111010101110111011001110011011101110111011100100111011101110010011101010011011101110010001001110001001001010111001000100111011101000111011101000011011001100000011101110111011100000111001000000111011101110010011101110000011100110111011001110111011101110111011100110111011101110101011100110101001001110111011101110111001000000111001101110111001001100111011101110100010101100101001001110111011101110111010100000111010001110111011100110101011101110111000001110111",
		"01110000001101110111010001000111011100110111011001110000000101010011001001110000010101100001011101110111011101100011011100010111011100110111011101110010011101110111011101110111011101110010000101000011011101110111000000110001011101110111011101110110011100100110011101110101011100010111011101100111011000110011011101110111011101110111011101110101010101100110011101110101011101110110000001100010000100100110011101110111011001110111011101110001011101110101011100110111000001110001011101110001010100110101011101110111",
		"01100101011101110111011101110010011101110111011101100111011101010011011100010011011101110111011001100001000000000111011101110101010001110111011101110100010001110111000101110111001001110111010101110011011100010000001101110111011101110101011101100111001001110011011101110110001000000111011101110001001100110111011101110100010001110011010100100111001001110111011101110010011101000000011000010101011101110000010101000111011101110111011101110010000101110111000101110000011101110100011101110011000000100011011101110111",
		"01000111011101110111011101000011011101100111001101110111010000010111000000100111010100110000011101000111011101010011010101000111011101000111011101100101011101110111011101110011000100010111010001000111001000010100011101110111011101110111000100000111011101110111010001110111011000110111011100100010000101010111011101000100001000100111001000100111011101110111011101010110001001110111011101110111001101110100001000110010000101100111011101110111001100110001000001110111001101100111010101100111010101110111011100100111",
		"01110001001101110100011101110111001001110111011001110111000101110011001001110111011101110111011101110011011001110111011101110100000101110111011101110101001100100111011101110111011101100111011101110100011101010111000000010111011101100001011100000111011101110111011101100111001001110010011100100101011101100111011101100110011101110000001000010111000101110111011101000001011100110101011001110111011000110111000101010111011101110000011101110010011100000111011101100100011100110111011000100111011101100111011101110110",
		"01100111001000010110001101110111011101110110011100000111011101110111000101110111010001000111000101110101011101010111010001000110011001110110011101010000011101110111011101100111011101110111011100000111011100110010011101110111011001110100000000010100011001100111011100010111011101100111011001110111001101110111011000110111010101110111011101110111001101110100011101110111011101010100001101110001011000010111011101010111011101110111001000100011011101010111001001110111001101000101011100110111011101110010011101110111",
		"00110001011101110111011101110111011101110111011100010011011101110111011100100100011000110111001001110111011100100111000001100111001000010100011100010111001001110111011101000111011101110000011100000111001001110011000001100111011101010111000101110111000101110111011101010010011101110111010100100010011100010111010001110111011100000000011101110111011100000111001101110111001001110111011101110010000001110111011100100001010001110001001001110111001001110011011101110111011100000110011101110111011100010111011101110011",
		"01110111000000010111011101110111011101110110011101110010000101110111001101110111011101110010000001000111011101110111011101110110001000110111000001110111001001110111011100010111011101110101011100110111001101110111011101110010011101110111011101110111011100100111011101110111011001100110011100100111011101110001011101110010011100010100011101110111011101110111010001110111011101110000011001110111001101110011010001110110011101000111011101110111000101110101011000110111001101110001001101110111001001110010000101110111",
		"00100111011101010101010101110111011101110111011100100001000001110101001101110111011101110010001001000111011101110101011101010011011101110100000101110111011100010111011101110111011100110111011101110110010001010111011101110111011101110111011101110111011100000111000001110100001100000111000000100010000101110000011001110011011101110011000101100111010101110111011101110110011101110001011101100001011101010011001100110111011101000010011100110000011001000011011101110111011101110111000001110111010001110110001000110010",
		"01110111011101110111000101110000001101010111001100110111010101110111011001110111010101110101011101110011001101010111011101110111001101110101010001110111010001110111010001110110011101110111011101100000011001110111001100110111000000000111011101110001011101100101000100110111011101100111011101110111011100100011011101110111011100000001010000110111000100110001011101110101000101100111011101100111010001110111011100010000011101110111001001110111001001110111011100010111011101110110000001110101000000010111001001000000",
		"01000111000101110111010101100000011100000111011101110111010001100111011101010010001001110111011101110101011100110111010101110001011101110011010100000000011101110000011101110100011100010111001101110101000101000111011101110111011000110001011101110100000001110000011101110001001001110101011100100111010101110111001101110111010001000110011100000111001001110111000101110111000001110111000101110101011101100111011101000111001101110111011101010111011100010111011000110000011100010111001100110111011101000100010101110111",
		"01110111011101000111011101110011011101110111011100000111011101110111000001010101011101010110011101110111000000000111001101000111011101110111011101110111001101110111010101010001001101110101011101110110011001110011010000110111010101010010001000010010011101000101011100010111000101110011011101110010010001110111010100010111011100000010011101110010000001110111011100100011011101110111001101110111011101110100011101110111000100110111001001110111011101110111011000000001011101110010010001110011001000110100000101010111",
		"00100111000101110111010101110111010101110111011101110111011101010111000101000111001000100111010001110111011100110111000000100100000001110101011101110111011100110111000001000111011100010011010101110111011101110000011001110011011101110111001101100111001100000111011101110111001101110111001101110011011101000111011101110111011101110010011100100100011100110111000101110001001001110111000001110111001000100010010000100111011101110100011100010111011101110010001001110111001100000101011101110111011100000111011101100111",
		"01110110011100100001011101000001010100010011011101110111000100100110011101110111011100010111011101110111011101110111011101010111011101110111011101110011011101110110011101010111011101110100000000000000011101110101011101110111001001110111000001010110011001010111011101110111001001110111010101110111011001110110011101110011001001100111011101110011011100100111001101110100010001110100011101110010011101110111011001000111010101110010011101000100001000010111011101110101000001110111001100100111011101110111011101110111",
		"01110010000001110101011100100111000001010100011000000011011100010000011101110011011100010111011101000001010001110100011101110001011101110111001000100111000101110101010101110110000101110111010101110111011101110100011101110110000101110111011101110111001001110111011101100010001101110011001001110111001100100111011101110111010001110101011101110111011101110111000101110111011101110010011101110111011101000110000100110111011101110111011101000111011101110011011101110100000101110111011101010111011101000111011101000111",
		"00110101001001110001011001110111011001110101011101110000000101110111000000110111011101110111011101110111000101110111001100000111000101010111000101110111010000000111001001110111011101110111011001110111011101110001011101100011011101110111001101000111011101000110011101000111000001110111011101110111011100010111011001000100011101110001011101010111011101110111011101110111010001000111011101110111001100100111001100010101011101110011011101110011011101110110011101110100011100100111011001000111011101110111010001110011",
		"01110001011100010111010001100111011101110111011100000111001101110011010001110010011100010100011001000111011101110100010000010111000101010010010101110101001001110111011101110111011100100011000001110111011101110111001001110111011101110100011101110100011101010010000001110111010001110000011101100011011101110110011101100000010101110100011000100101011101110111011101100001001101110111011101110010011101000001010001110101011101110111010001110111011101010111010001000111011101110010011101110111010001100000011101110111",
		"00100111011101110111001000110011011100100111000100000111000001110111000001110111011101110011011101110101011101100111001101110000001101110111011101110001010001110111001001110110011100110111011001110011010000010110011001110010011101000100001100110111011101110111011101110111011101010010001101110001011001110111011000000111001001010101011101110111011001110111011101110111011101000110011101110110011001000111011101110101011100000011011101010111011101110101011101110111011100100000011101110111011101110110011101110111",
		"01000111011101110111011101110001011101110111000101000111011101110111011101110111011100000111011101110000011101110111011001110110010001110110001100010101000001110001001001110111011100100000011101010111011100100111000001110111011100100110001100010101011101110001011101110001011000110111011100100101000001000010011101110111000000010111000100100111011101110101011101100100011100100111011101110000011100000111011101110111011100000000010001110111000101110111001101110111010101110000010001110000011101000000011101110000",
		"00110101011101110111001101110111010000110100011101100111011100110111010101110111011100110111010100110100011100000111000101110111000101110110000001100111011101110101011100000111011101110000011100000100011100100111011101110111011001110111001101010001011100110111011101110111011101110111001001110111011100010011011001110111001100100111011100110010000001110010011101110111011101110111001101110111011101110111011101000111011101110101001100000111011101110111000001110101010001110111011101000011001101110000000001110001",
		"01110111011101000111000101110000011101000111011100010001011101110111000101110010010001110111001101110011011100110111011000100111011101010010011101110110011101110110000101110111010101100000011101110100011101110111011101110111011101000111011100100100011101000001011101110000000101110101011101110111011101010010000100010111011101110011001001100111010100100010010000000111010001110111011101110110011101110111010001110110010001110111011101110111011101110110011101110110011101110111000001010111011100010111011101110111",
		"01110000011101110010011101110111011101110101011101110011010000000110011101110111011100100111011101110101000000000111001001110111010100100100011100000110001101110111011000100111011101110111000001110111011101110111010000100010011100110000011101010101011101110000001001000111000101110010011101110111011101110100011101110011010001110111010101110010011101110111011100000001000101100010011101110000011101010101011101010111011101010111011101000101011101110111011100110110001101110111010101110111011001110001011101010011",
		"01110111011100000111011101110010011001110111011100110100011100010011011101110111011101110111000001110100010101110111001000100001000001110110000001110000000000110000011001110001001101110000011100010010011000100011000101010100011101110010001101110010011101000001000101110110001101110111011101110111011101110010011101110111001101110101001101110100000100110111011100110101011100000111011101110010011101110111011101010111011101110000011101110111010101110110010100010111000000100011010100110110011100110111011101110101",
		"01110101000001110111011101110111011101110100011101110111001001110010011101110101010101000111011101110111011100010111011101110111001100000010011101110011000001110011001101110000010001010010011101010011011101010000011101110110001100010100001001110111011101110111010000100000011100100111010100000111011101110010000001110111011101110111000001110001011100010111001001110110001101110101010101110110011101000111001001110111011001110001001001110111011101110000011101110111011101110001000000100111011100100111001101010110",
		"01000111010101100111001101110111000100110111011101110111011101110111011101000111011001110101011101110010001001110111011001110111011100110010011101110111011001110101011101110110010000010100011101110111011100000111011000100011001000010111000001110111000101110111011100110111001001100111001101110111011101110111000000000001001000000111011101110111011101010001011101110011010001100101001001110111000101010111011101110111011101010100001100010001011100110010010001110101011101100111000101110111011101110110011001000010",
		"01110111011101110010011101110111001000010100000101110101011101110111011101000111011000010111011100110011010001110001010101110111011101110101010000000111000000010101011101100111010001110111011000010111011101110110011101110111011101110111011101010111011101110110001001110111001001110111010101110010010001010100011100000011010101110000011100110111011001110111011101110111001001000011011101110111011001110000011000000111011101000111000001110111011101110000011101000100001001110111010001000000011100110000011101010001",
		"01110111010001110111001000010111011101110111011101110111001100010111011000110111011101110000000001110100011101110111000001000111011101010100011101110111011101110111011101110100011100010101011101100100010001110111011101110111011001110111011101110111011101110111011101110111010101010011001100100110010100110111000001010111011101110111001000010111011100100100000001110111001101000111001001110111011101110110010101110111010001110111011101110001010001110111000101110101000101110101001101110001011100000100011101110111",
		"00010010011101110001010101110101000001110100011101110111011101010111010000100111010001110111011101110111011001110101011101110000011101110010000000110100011101110111011101110111011101010111010101110111010101110111010101100111011101110001011101110111011101010001001101100111011101110011011001110111011101110001011100010010011101110101011101010111011100010111010101110100011101110001000101110111011101110110010101110111011001110111000000110111000101110001011100110100011101110111011001000100000101100111011101110111",
		"01110100011101110111011100110111011101110111011101110111000101110101011100010101001001110000011101110111011101110111001101110101001101110111000101110111011100100111011101110111000001110111011100000111011101110111001101110000011101110111001001110110011101100000011101110101010001110011011100100000011101110111011101110111011101110111010001000111011101110111011100100100010001110111011101110111011101110000011101110111011000110111011001010111010100010000001000100111011101110111011101100100011100100111001100110111",
		"01110111011100000100011101110111011001110010000001110001011101110100011001110110010000100101010101110111011101110010011101110111011101110111010001110111000000010111011101110111010000110100011101110001011101110111010101110111011101110110011100100010001101010000011100000111011101110110011101110000000001110111011001100111010000010111011101110111010101110101011100110111011101110111001000100000011100010110000000110111011101110011011100010101001100000111000001110111011100000111011100100111011101110111011101110011",
		"01110111011100110111000101110100011101110111001101110000011101010111010001110111010001110000011101110111000101110000011101110111000101110111000001010111011101110011010000110110010001110111011101110111000100100111011101100111011100010111011101010011011101010111011101000111011101100100000101110111010001110101011101110111011101010000011101110010011101110111000101100111010000100111011100100100010001110111011101110110011101000100011101100100001000100111001101110010011101110111001001110111010001110001011101110111",
		"01110011010000000110011101110110011100110111000100100111010101110000011001100001010001110010011101110111011101010011011101110111010101110111011101110100011101110010000001110010010001010111011101110111011101110111011101110100011101000111001001110000011100110011011101110100001001110111011101110111001001010100011101110011001001110111001000000011011101110111000100100010000001100111000000110101011101110101010100110111001101110110011100010110010100100111010001010111010101110011011101110010011100100111001100010100",
		"01110001010000010111010101110110011101110111011100010000011101110111011101110111011101110111011101010111001001110010011101110100011101110010001100100111011100010001011101110111001101110001011001110001011101110111011101110111011101110111011101110101000101110000011100000011011001110101011101110111001001110111010001110000010100110111011001110111011101010111000000110111011100010111011101110111011101110111011101100111011100010100001001110111011100000000011101110010011101110111011101110111000101110111000001010111",
		"01110111011101110111011101110110000101110111011101110111011101110011011101100110011100100111001001110111011001110010011101110000011101100001001101010100011101010010011101100111001001110111011101000100011000100001000000110001001001000000001001110000011101110101011101000111011101110111011101110111010101110011011101110101000101110001011101110111011100000111011101110111011101110000000001000110011101110111011101110111000101110111011101110011010001110111001000010111010001000001010101110101011101110111011101110111",
		"00100101011101100011010001110111011101010000011101110111011100110111001001110111011100100111011101110111011001110101011101110111010001110110010000010110010101110100011001110111011101110001011101110101011000000011011001110111011101100111011100000110011101110101011100000111010101100111011001010011001101110100011101110110011100010011000101110011000001010100010000000011011100110011011101110000011101110111001101010111011100100011011101110111011101110111010001110000001001010100010101110111000100000111011101110111",
		"01110011011100000100011001110111011100110111011100100111011100110110011101110010011101010000011101000000001100110000011101110101011001100101011101110111010101110111010001110001001101110111011100100111011101110111011100110111000001110100001101110100011100110111001001110101000101110101001101110101001001110111011100100001001000100111001101010001010001110111001001110100011101110110010101110111011101000111011101110101000101110111011100000111010101100111011101000001001000000111011001010111011101000111001101110111",
		"01000111001001110111010001100100011101110010010101110101011101110001011101110111000001110111011101110111000100010111011001110000011101110010011101110111011101110111011100100101010000000111001101110111011101100111011100100101011001110111011101110111011101110111011101110100011101100001011101110001011101000100010100000010011101110001001001110111001001000100011101110111010001010111011101110110001101110111000001000111011101010111011101100111001100000111010101110111001101100110011001110111011101110111001101110111",
		"00010101001101110111011101010101011100010111011101110111001101100111011001110111000000110010001001110010011001010111011101000111011101110100000101010111011101000101011001100001011101100111001001110111011101110100001100010111010000000111000100100111011100110111011101000111001001110111010001110110000101110111011100100101011101110111001001110111001101110111011101110111001101000111001101110111010101110000011101110111011101110111011101110010010001000011011101110010001101110110011101000101011000100110010101100111",
		"01110101011101110111000001110111001100100111011101110111011101010101010101110111011101110111011101110001011101110111010000100010011101100111011101000111011100010111001001110111011101110111011101110100011101110111010001110111011100110100000101110110010100010111001101110111011101110110011000010111011101100000010101010010011101110111001001110111011101110000011100100010011101110111011101110111011001110111011001110111011101110001000001110111001101110111011100110111001000010010000000110011011100000011011101110111",
		"01100111001001010111001101110101011000010111011101110111011101110111011101110111011001000111000101110011011101110111011100110111011101110111011100110111000000010100011101110111001100010111011000110111011101110100011101110110011100100111011101110111011101100111011001010111011101110111010001000111010100110010000101110001011101110111011101110111011101000110011101110000000001110011011101000111011100110111011100010111000001110001010001110111010101110010011101110101011101110111011100010111011101110011011001110101",
		"00000111011101110111010001110111011101110111011101110111000000010111001101110111001100100101011000110111011101110111011101110111011101110001011100110110010001110111011100100011011101110111000100100110011101110000001001100111011100010111011101110111001001110111010001110111011101110110011101110111011001110111010001110111011101110111010001110111000101110101010001110111011100110111011101110001001101110111010001110111000101110000011001000111011101110111011101000111001101110111011101110000011101110111011101110111",
		"00110100011101110111011101110011011101010111011100000101011101110111000101110111011100110111011001110111011101010111010000100100011101100101011101110000011101000111011101110111001001010111011001110111001100100111011101000101011101110111010101110100011101110010001101110111000001110111011101100011001001110010011101000111001001000111000001110010011101110101011101110110001101110000010001110111011101110111011101110010011101110111001001110111011100110000011101110011011100000011011100110111011101110111011100010001",
		"01110111001101110010011101110111001001110111000001110011011101110111011101110111011001110111011100010111010001000111011100000100001101110000011100100111001000010111011101110111001001100011011100000111011101110111011101110111011101110100011100110000000001010111011101110111001100000111000001110111011101010100011101010001010101110011011101110111001101010111001001110011000000110111010101110001011100010111001001000110011101110111011101100000011101110111011101110111010000000111011100010000011000110111011101010111",
		"01100010011100110111000101110111011101110011011100100000011101110110000101110010010101110111001101010111011100000111001000010110011100010111011100110111011100010111011101110000011101110001000000110111011001110111010101110001011101110011011101110111001001000111001101110111011101100111011100110111000001110111001000000111011101100110011100010101001001110111011101110111000101010101011101110111011101010110011101110111011101110111011100010111001101110111011000110001000001110111011101110111011100110000011101110111",
		"01110110011100010111011101110101011101110111011100100111011101110110010101110000011101110001011101110111011001010111001101110111011101110101000101110111011101110001011001110101011101110111010101110111011101110111011101110111001101110110011101110110000101000011011100000101011101100000011101110111000101010111000001110010000001110010011101110111011101000111001101110111011100000111011101010111000101010010011101010110010000000101011100110111011101000000010101110111001100110111001101110111011100100111010101110111",
		"01110001011001110100011101110111011101110011011001100111010000100111011101100111000000000111001000010001011101110000011100000000011101110111011101110011011100100111000101110110011100110110011101110111011101000011010100110111011101110111001001110111011000110101000000000111011100000111000101000010011001010100011101110101011101110110011101110111011101000111010001010111001001000111001001110111011100110111010001110111011101000101010101110000011101110111011101100000000001000001011100000111011100000111000101110100",
		"01110011001101110110010000010111011101110111011101110101000001100111011101110010001000010100011100000100011101000001011101010111000001110111000001010111011100110111010100010100011101110100011000100111011101110110011101110111010001110111011101110010001001110111011101110111010001010110011101100011011101110000000001010010011100110111011100010100011100010000011101110111010001110111001101100111011101110111011101010111011101010000011101110011011101110011011101110111011100000111001101110111011001110111011101110111",
		"01110111011101110111010001110111011101110111000001110010010000110111011100110010011101110010011101110110010101110000011101110100011101110001000001110111001001110111011101110111010001110111011100110111011101110111011101010010010101110010011101110111011101000110001001110111011101100111000101110111010000010011011101110111011101000001011101110111000000100101011101100011010001000100011101110111000001100111011001110111011101110111010001110111001000000111011001110111011001110011011101110110001100010010011100100111",
		"01110111010001110111011101110111010100100111010101110100011101110111011101110111001100100010011100010111010000010001011101110100011101110111000001100111001000100101011100000110011101110111011101110000001101100111001000100001010101100000011101110111011101110101011100110001011101110111010101110111011100100000011101110000001001110111011101110011011101110111010101010010011001100111011100100111011101110000011101110111011101110111011101010111011100110001001100110000000000100111011101000111000001110111011101110111",
		"01110111001101110111011101000001011101110111001101110101011100110111011101110010011101110011011001000111010100110111011100110111011100000011000101110111000001110111011001110111011101010000011101100111000001110011011101110111011101110111011101110111001001110000011101100111011101100010011101000011001101110111001101110111011101110111000101100011001001110111011100000111001101110110010101110111011101110011000101000110000100110111011101010111011001000101011101000000011101110111011101110111011101110111010001110111",
		"01110111001101110111000101110000011100000001011101110111010101110110011000110111011101110111010000010000011101000111011101110111011100000111011101110111011100110000011101100111000100000111011101110000011101010100010001110000000001110111010001110111000001110111001000000110011000000111011001110000011101110111001101110111010001110101011101010000001100110111011100000000011101110111011101110001011001110111001001010011000001110111011100000000010001110111011101110111011101110111001101110111000100010001001100010111",
		"00000111011101110111001101110111001101110111011100010111000000110010010001100111011101110111001101110011010101110111000101110111000000000111011101000111011100110111011100000101011101010100000101010111000100000111011100000111011101110111011100110111011101100111011101110111011101100111001001110111010101110101001001110111011101110011011100110111010100100111010001110111000000010110011101110111011101110111011001110000001100000111011101110111001101110100011001110111011101110111011101110000001001110001011101110111",
		"01110101011101110111011101000011011101110000011101100111011101110101011101110011000101110111011100010111000001110111011100010111000000100101011100100100011101010100001000100010010101110111011101110111001101110001011101010111001101110000011101110111011101110111011101000111011101110111011001110111010001110111010100110010011101010001010101110011011100000011001101110111000001110111011101110111011101110110010100010111001001110111011101110111000001000110010000000111001001110111010101110111011101110111011101110010",
		"00100010010000000000011101110101001101110101011101110000011101110111011101110111011101000110011001000111010001110111011101110011011101110111011101110000011100100111001101110111011100010111011001110111011101110111011100100111011101110111001000100111011100000111011101110111011101110111011101110010011101110111001101100111011101110000011100000111011101110011001101110111011101110000001100010111011100110101011100100010011100000100001001110111011100010001001001110111011101110100000101110111011101010110000100100111",
		"01110111011100010100001100100111011101100111011101110100000101110111000101110111000001100000001000100000011101000101010101100100011001110111000101000011000100010111011101110111011001110111011101110111011100000111010001100111011100010111010000010110010001100010011101110111011100110111011000100101011100110011000001110111011101110111011101110111001101000010011101110110001101110111001101110111011101110111011101010111000001100111000100000100001000010111011101000111011101110010011101110111000000110111011101110111",
		"01110101000001110010000101110111011100010011010101110111010101110111011101110111011101010111011101110111011100000101000001110011011100000011011101110111011100110110011001000111001100100110011100100111011101110001011101110111001001110011011100000111001000110110001001110111011101110001000101110111011101110111011101110111001100100101001101110111001101110111011101110101011101110111010000110101011101100011011101110010000101110111010101110001011101110111001101000000000101010001011100100111011101010111011101110111",
		"01110111010101110111011000100111011001110101001101100111001001110101011100010110011101110010011100010111001001110000011100100111011101110111011101000111001001110111010001110111001001110110011101110111000001110000000001110111010100010111001101110000011100010010011001100111000101000111010000010111001101010111011100000111011101110111011101110010011101010110011101110111000001110101001001110010011101110111000000010111010101110111011101110010011101010000011100000010011101110000011101110111011101110111001000000111",
		"01110101001100010110000001000111011100110111010100100010011001110001011001110111011000100101000001110110011101110111011101110100011100010101011101110111011101110011011101110100010101110100011101110111001000010111000101110111011101110111001001110100001101110010011101110001000001100101011101110111001001110110011101110000010001110001000001110110000101110100011100010101011101110010010101010111011101110111011100100110011101110111000001110111011101110110011101110111000000000111001000110000010000100001000101110111",
		"01100110011101000001011101110100011101110111001001110111011101110111001000000111011101110111000001110111011101110011011100100101011100110111010101000111011101110111011100010111011101110111011101110100000101110000011101110010010001110011011001110100011101000111011101110111010001110111011101110011001001110111011101110011000101110101011101110111011101110010011101000001011101100111011101010000011101110111000001110111011100100001011001100111010101100101011101100111011101110111011101110111000101110111011101110111",
		"01110000011101010010001001110000011101000111011100110111011101110101011101000010000001110111011101000111011001000100011100000111010001110111001101110111011101110101011101010000011101110111011001110000010101110111011101110101011101110111011101110111011101010111000000010111011101000111001001110111011101110110011101110000000000010111000000010100010001110000011101110011011101110111010101110110000101010111001101110101011001110111011101110111000101110010000001110001000001010101011100000010000000010001011101110111",
		"01000110000000010111011100110111011101110111011101110111001101110010000100110111011101110111011100110111011100100001010001000110001101110111011001110111000100010110011101110111011100010111010101100111011101110111011101110111011100010010011100000111011101110111011000000010011101100100011101010111011101010111010001000111011101110111000101110111011100010010011101110010011101010010011100000111011101110100011101110011000101110110011001110001011101110001011101110111011001110111011101000111010101110111010001110111",
		"01110111001000100111011101110111001000000011010101110111001100100111011100000011010101110111001101110111000100100111000100100111011101110111011100000101011101110010011101110111000001110111010101110001011101010001011101110001010001110111011101100110011101110111011100010111001001100010010101110111011100000000010100000011001001110111010101110110000001110111011101000111011101110000011100100111001001010111011100110111011001100111001101110100001001110111001101110111000101010011010001110011011101110111011101110000",
		"01010111001100100111001100110111010101110111001001010111001101110010011101110010011100010001001100100001010001110010011100110100000100100011011101000111011101000111000101110110011101110111011101110011010001110111011101110111001001110111011101110111001001010111011100110111011101110001011101110011000000010111000001110101011101110001011001110011010101110111011101110001011101110111010101110001011101000111010101010111011101110101011101110001011100000011011101110111010100100000011100100001000101010111011101110100",
		"00100111011101110111000100100111011101110111011101110111000000110000001101110011000001110111010001110111000001010010011000100110011101110101001001110001001100100111010001110111011101110101001101110111011101010100011101110111011101110001010101010111000000100111011001000100001101010000011101110111011101110011011100010111011101110111011100010110011101110111011100100111011100000111011101000111011001110111000000010101011101110111011101010111011100000011010001000111011101110101011100100111011101100111000101110111",
		"00100101001100000111011001110111011101110010000100110100011100000111011101010111010001110111011000010111011101000100011101110100010101110101011100100011011001110111011101110111000001110111000101110111011101110101000101110000001001110011011101110111011101000111011101100111011101110111011100110010010001000111011101110001011101110010011100110111011100100101000100010111011101110111011101110111000100100111011001110111001001100111000100100110010001110111011101110010011100100111000101010111011101110010011100100101",
		"00010111001000110000010001110111011101110111000101100011000101110111011100010000010001110100010001110001000001110000011001010111011101000001011100100000001100110111011101010101001001110111011101110111010001110111011100110111011101110111011101110111011100110011011101110111011101110011010000010110000001110111001001110111010001110111011100010000001101110011000001110111011100010000011101110111011101110110011101000000011101110101011101110111011101010110010101110101011101000111010001110111011101110010001101110111",
		"01110111011100010111011100110111011101110111011101110110011101000000001100000000010000100010000101000000011101110000011101010001000101110001011101110000000000000000011101110111011101110100011101000100011101110111011101110111011101100011011101110111011001110011001000110000000101110001011100100111011100100111010101110111011100100111011101110101011000010111011101110110011100100011001100000111011101110110011101110011011101110111001000000111011101110000011101010110001101110111011101000111011100110011000101110111",
		"00100111011100100100000100100111011101110111001000000111011000010111001000010100000000100111011101110111010001000001011001110111011100000110001101110111001000010111011100010111011101010111001001110011011100010111001001000110011101110111011101000111001100000111001100010000001001000011010001110111011101110111011101110110011101000001011101110100000000010111000001010011010100110111011101110111010101110111011100110110011101110111001101010111011101110111011100100111010101110111001001000001011000110111011101110100",
		"01100111010101110000011101110011010100000111001101000111001101010111001101110111011101110101011101110001000100000111011101000111011100010111011101110101010001110111011101110010011100100101011100010110011101110011011101110010011101100111011101110001011101110111011100110101011100100110011101110111011101110111001100100111011100100001011100100110010101110110011101000011011101110011011101110011001001010111011101110010011100010111001000000001000101110111001101110111011001100000011101110111011100000110011101010111",
		"01110111011100010011011001110111000001000001001101110111011101110111011101110010011101110111011001110111001101000111011101110001011101110100011101010111011101110011011100100001011101110111011101100101011101110111010001110111011101110010000101110111011001010111010001000011011100110111011001110111011100100100011001000111011001100011011101100111011101110010011101110111001101110111011100100111000101110111011100100010000001110111011101110100000001110010011100010111011101110111011001110111010101110111011000110111",
		"01110111011101110010011101110111001101010101001001110110000101000001000001110111001101110111010001100111000101110111011100000000000001110111000100010111001001110000011101110100011101010001011001010010011101110111011001110000000101000101010101010111011101110111011101000111011101010111011100100001010000000100011101110111000100100111011100110101011101110111011100010111011100000110000100110111011101000111011001010111011101000011011101110111000000000111011101000111010001110111000101110000001001100111010001110111",
		"01000111001001110011011100010011010101110101011101110111011000000011011101110111010001110111011101110101000101110111000001010111000101110111010101110011011101110000011100010001000001110100010001000111011100110111001101110111000001110011011101110101010001000001011101100111010001110110011101110111011101110101010000110111000001000111011100010110011101110001000101110111000001010111000101000111011101110100000101110111011001110111011101110111010000010111010101110001011101110011000001110001011101000010000100100111",
		"01110111011101000111011101110101000100010111010101110110011100110000011100100111001100010011011100100101001001110111011101110111000001110000011101110111011101110111011101110111011101110111011101000111011100100111011101110110011101110111011101110111011101110111010101110111000000010111011101110111010001110100011100100111010001110111000101000001011101110100010001010111011001010111011101110111011101100111011101110001001001100110011101110111011101010001000101110000000000000111001000000111011000110111011101110111",
		"00000000011101110111011101010111011101110100011101110111010000110100010101110111011101110011001101000111011101110111010001110111011100110111001001110111000001100000001100000111011101110110011001110011011001000111011001110101011101010111011100010111000000000111011101110111011101110111011101110111011100100000000001110101010101110111011101110101011101110010011101110111011100010111011101110101000001110111000101110111001101110111011101100111011100110111000100000010011101110001011000100010010101000011011000000110",
		"01110100000000100111001101110000011101000111001100000111011100100111011101010111011100110101001001000111011101010010011100110100011101010111011100010010000101110001010101110111011101110000010101010111011101110111010101110111011101110111000100100111011101110011010001000111011100010111011101110111011101110011011101010111001101010111011100010000000001110110011101010111011101110000000000010111011100110111011101110111011101110001011100100111011101110000000001110111011100100101011101110111011101000011011100110111",
		"01110001011101110111001101000111011100000111010001110100011100100111001001110111011100000001001001110101011100110111011101110001000001000111011101100111001100010111011101110011011101110000010101110000010101010111011101110111011101110111011101110111011101110010001001110111000001100111001001110111010000100111010001100010011100010111011100010111000000000010011101110111011101110111001100010111011101110000011101110111000101110011001101110011011100010111010001110111000000000000011100110111001001110111011001110111",
		"01110111011100010001011101000000011101010111011101000010001101110111011101110111000000110011011001110010011101100111011100010010011100010000011100010111011100110001011101100001011100010111011101110111011100000111011100010100000101110111001101110111010101100000011100000111011101110111011100100111011101000111010101010111001001110111011101110110001101110101010000110111001001110111010001110001011001110010011101010100000000000111001001110111011100000111011101000001011100010000000101000001011001110111011101000111",
		"01110111011101110111010001110100011101110110011101000110010001010111011101110111010001110111011101000111011101110111011101110111011101110010001101110000011101110101001101000101011101100101001101110001011101000111011101110110011101110000001000100100001001110111001001110001011100110111010001110111011100110111011100010101000001110001001100000000011101110111011101110111011101110111011100000111000100100111010001100111011100000111011101110110011101100001010101000111011101110101000100100111011100100100000101110000",
		"01110111000100100111011100100111010000110110011101110101001100100111000000110000011101110101011101110111011100010010011001110000011000100111011101110111001101000111011101110010011101010010000000100111011101110011010000100111001000000111011101110000010101110101011100100011011100100111001101110111011101110111000000010010011100110101000001000100011100100111011101110100010101000111011001110111011101110100011001110111011101110111011100000001001100010111011000100111011101110110011100110111011101110111011101110111",
		"01110111011100100111010001110000011101110110011101000101011100010111001101110111000101010111010101110111011100100100011101010111011100110100001101110101001100100111000001110111011101000111011100010111011101110001011101110111011101110010001101110100011101110111001001110111011101000111011101000010011101110111011101000111011101110111001101110011001101010110011101110100011101100111001001110111011101110111011101110111011101110000011101100111010101110111011101000111011101100101011000110111000001110111000001010000",
		"01110111001100100111011101110011011001110101011101110000001101110111011001110111011101100111000100110111011100000000011101110110001101110111001101110111001101100111011101110111001101110100011101110111011101110110011100100000011101110111001001110111011101110110011101110100011101110001011101110000011100000111011100000011001101110111010101110111011101110111011101100111010100110111011101110111011101110111000101110000011101010101011100110101011101110111010101110101011001100111010101110110001100110111011100100001",
		"00100111011101110101011101110111011100010111011101110111010100110111010001110111011101110100011100110111000001100111011100010111011100000111011000000111001100010111011101110111011101110001010000000111011101000111000001110101011101110111011101010010011101100111011000100011011101110001001101110111010001110010001101110001011100000111011101110111000101000111000001100111011000010111011101100011011101010111011100000111001001100111011101000001010001110010011100110111011101110000010101110001010001110000011101110111",
		"01010111011101010111011101110000011101110100010101110111001001110000000101100101011101010111011101110111011101110111011100100111011000100001011101110100000101110111011100000111010001000001000101110111010101110111011101110010001001110111001101110111011101110111010000100111011101000111011101110111011100100111001001000111011101110111011001110100011101100111010101110111011101110110010001110110001101110100011101110000011101000111011101110111010001110011000001110010011101110111011101110111011101110111010001110100",
		"01000111011100110111011101110111010101110110001001110111000101110000011101110101011100010010000100100111011101110111011101110111011100110001011100010010011101110111011101110010000001110111011000000111011101110111011101110111011101110010000001110111011101000111011101110111011001010100011101100100011101010111001101110011011100000111011100100110010101000110000100010111010101100100001100010011011101000111011101110111011101100001011100100111011100110111011101110010011001110111000000100111011100110000011101010111",
		"00010111000100100111011101110010000100110111011101010001011101110010011101110111011101110110000101100001011101110111011101000111011101110111010101110111011101110111011101110111010101110110011101110111011101110111011101110111011001110111011100000010011100100010011101110111000101110111010101010000011101110111010100110111001100100101000001110111011100110111011101110100011101110100011101110011010101110000011101110111011101100111011101010111011101110111010001110111010001110101011101110111011101110000000101110011",
		"01010010001100000111011100110101011100010110011101000111001000000101011101100111011101110111011001110111011101110100011100100100011100100111011100010111011101110100011101110100010101110000011101110100011001110010000001110111001000100001011100000111001001110010000000000110011001000111010000110111011101000111000001110111011101110111011101110111011101000111011100110100011101110101011101110111011100010111011101110000000001110111000101110111011100100111010001110111011100100111001001110000011101110100011101110111",
		"01000110011101110111001000010100001101110101011101110111000001110111010101110111001101110111011101110111011100100000011100110110011101110011011101110111011001110010001100110111011100110101000000110111011101100001010101110010011100100000000000100100011101110111001101110111010001110100000101010010011001000101011101110111010101110111011101000111000100100111011101010111000101100101011100100111011101110010011100100111010100000101011101110100011101110111000000100111001101110111010001110110011101110111011101110000",
		"00000010011101000111011101110111011001100111011101110111001101110111011101110100000000110111011101110111001101110111010000010101000000110000000101110111011100110010011101100111011101110111011100010111010101110111011101010010010001110111011101110110000001110111011101110001011101000110011001110111011101110111000000110010000101010100011101110110000101110101011100100111011101110101011100100111001001110111011100000100011101010111011101010111011101110111011101110111001101110111010100010111010101110000011101110101",
		"01110101011101110111011101110111011101110110001100100100011101010111011101110110010101110011011101110101011101000001011101110111011101100111011101110111011001110111011101110111001001010101011101110111010101110101011101110100001000010111011101110100011101110111011100010111001001110011011101110111011101110111000101110001001101110101011101100111000101110101001001110011011101110111011100000111011100110111000101110100010100010111010101010111001001110111010101110110010001110110011101110110000000010011011101000111",
		"01110111011001110011011101110111000000010111000001110110001001110111011101110110011100110111001001110111011101110111011100110111011100100111011101110111011100010101011101000111001101110100000101110100011100010111010101110111011100110111011100110111011100100010000001110011000101110111000101110111010101110010011101110111011101000111001100110111011100010111011101110111010001110111011101110110011101110111011101110111011101010010000000100100011100010111011100000110011100110111010001110111011100100001000101110011",
		"01110111010001110111001001110111011101000111000001110111011101110111011101100111010001000011011100100111011101100111011101110111010101110111010001110111011101110110011101110110000101110111010001110001001101110111011101110111011101110111010101110111011100100111011100100111011101110111011101010011011101110111011000010001010001110111010101110000011101110000011101110101011101110110001100100111011101110111000000000011011101110011011101110001011101110111011101010100011101110111011101110111011101110110010100000111",
		"01110111011101110111011101110111000001000111011100000111011101110111011001010011011101110111011101100111011101100110011101110111010101110111000101110010011001010111011100010111011001110101000101110100011100110111011101110111001101110000011101110111011101110001010100010111011101100111011101110111010001110101011101110111011101110100011100000010011101110111000000010111000100010111011101010001000001110101011100100111011100000000011101010111010001110111011101110111011101010111011101010101011100100111011101110001",
		"01010111000001110110011101110111011101010111001001110111011001110001011101110011011101110110011101110000011101110000011101110111001101110111011101000000011101110111011101000010011101110001001001110100011101110111011101110111011001110111001101110000011101110011011101110110010101110000011100010111011101110111011101110111011101010000000100110111011101000111011101100110011101110001011101110111011101110011010001110100000101010101011101110111011101110000011101110111001001110111011001110111011101110111010001000111",
		"00110001011101110100001000100000011101110001000001110111011000100111011101110111011100010110011101110000010001110111011101110111011101000111011101110111010001110100001101110111000100000010011101110100001000100000010101000111011101110111011001110000011101110111010001000111011100100111000101100111001101110111011100100111011100010111000100010111011001110111011101110101011101110111010101110111010100110111011101000111010001000110011101110000011101110110011101110111011101110000011101110101010000100010001101000111",
		"01110110011101110111011001110101000100000111011101110001011101110111010100100010011101110110000100000111011100110111011101110111011101010110011101110111011100100111000101110011001000010010011101010000011101110111011101110111011101110111000101110010011101010111010100000101010100100111011001110001001101110111011101110110000000110001011101110100011000100110011100000111011101110111010001110000011101110111010101110111011101010111011101110111010101110111011001100111011101110111000101110111011100100101011101110110",
		"00000011011101100100011101100101011100010100011101110011010000100111011101100100011100010011011000100011011101110010011101110111011101100011011101000010011100000101011101100101011101110111000001110111011101000101011101100011011101110111000100000111011101110111011101100110010001110101011100100111011101010111011101110101011101110111011101110111011001110101011101110000000000100000000000100111011101010001011101110111010001010111011101000111011101010011011101110111011001000111011101010011011100110111000101100111",
		"00010111011101110101001000010111010000100100011001110111000001000111001001110111011100000000001101100100011101010100011101110011001101110001011101110110011101110111000000100010011000000111011101110111011101110111000001110100011100010110011101110111011101110011011101110011011101010111011101110000011101110101011101110101010001110100010001110111000101110000011101110111000101110111011101100111010000110111011101110111011100000100011101110111011101010110011100100111011101110111011101100111001101110111000101110110",
		"01010111010101010111011100010110011100110011000001110111011100100111011101010001000001110010001001110110010101110110001001110111011101110111011101010111011101110111010000110111000000000010011100010110001101110111011001110111011101010111011101110101001101110110000000000111011101110101011101000010011101100111010100010111000101010111001101110000000001110111011101110111011100010111001001110111001000010111011101110111011101110111011100000010000101110011000000010100001100000101000001110111001100110011011101110111",
		"01110101001001110011010101000001010001110011011100000101010101110011011101110111011101110000011101110111010000110111011100000111000101110111011101110011001001100111011101110010000001110100011101110101001100000111001001110110011101000101001101110110011101110111011101000111010101110110011100010110011101110111000001010111011101110010000000100111001001110111011101110111011101110111011100110000000101110111000101100111011001110101011100100010011100110111011100000011011101010001011101110001011101110111011101110000",
		"01110000011101110111011101110111011101000111011101110100011101110010010101110111010001110010011101100010010001110101010101000101011101110111010001110010011101110111010001110111011101110010010101100111011101110111011001110011011100000101010100100001000000100111001001110111011101100111011101110111010001110110011101110111001101110110010101110111011101100011011101110110011100110100011101110001011100110111011100000111011101110100011001010001011100100111011101110111001000110111000000100110001101010111001000010110",
		"01110110011101110110011101110111010101110000011101110000011101110111011001010000011101110111001100110111001101110111011101110011011101000111010101010010011100110111000001110111000101000111011100000011001001010111011100000110001101110000001101110111011101110001011100100111011101100111011101110110000101110010011001110111011101110111001001010000011100110011010101000111001101110111010100010111011101110100010001110110011101100111011100100100000001110111011101100111010101110111011100000111000001110111011101110111",
		"00110111011100100111001001110010011100000111011101110101000001110111011101110111011100010111011100010101011101110111001101010111011101110001011101110111011001000011011101110111011101100111011001110110011100110111000101110010001101010111000101110111011001110010000101110111011101110111011101110111011101110100001001110000011100110000011001110010011101000111011101100001011101010111001101110011001001110111011100100111011101110111011101010111011101110111011101110001011101110001011101110101001101110111011101110111",
		"01110101001100110001011101110111011101110111010001000100011101110111011100010111011101100101000100010111000100100111010101000000011101110111000101010111011101110010011101110100001101110011011100100011000001110001011101110111011101110001011100000010011100000010011101110111000001110101010101110111000101110100011100100010011101110111011100110111011101010000011101010000011101110010011101110111010001100111011100010111011101010111011100000111000100110111011101110001001101110001011101110111000001110110011101110111",
		"00000000011001110010011000110111001101110111000001110111010101110111001101010010000001000000001001110111000000110111011101110111011101110110010101110000011100000111011101110000000001110111001101000111011101100010011101110010011101110000010101110111011101000111011101110110001101100100011101000100011100010111010001110000010100000001010000010111011101110100011001110111000001110111001101110111010101010111011101110111011100000011000100110011011101010111011101010111001100010111011101110011011101110100011101110001",
		"01110000010000100111011101110111000001110111011101100111001000010111011101110111011100110111011101110111011101110001000001110111011101110010001100010111010100010001000101110111001101110010010101110111011101100011011101110111001101110111011101110111011101110111010000100011011101110111010100010001011101110111011101110111000101110100000100100111000000010111001001110111011101000111000000010111011101110111011100110011010001110111011100000100011001100111011100110111011101110111011101110111011101110000011100000110",
		"01110011011101110010011001110111011101110111000001110111001101110111011101110111000101010011011101110100011100010011000101110110001001110111011101110111011101000111011100100100011100100111011101010001001001110110001001110101001001110111000101010101001101110111011101110101000101110010000100110110011001110111000001110100011101110111011100010110011100100111011101000110000101110111011100110111001000010011001000010111011101010111001101100010001001110111011101110111011100000111001001110010001001110111010001110111",
		"01110011000101110110000001110111000101110100001000100010011101110111011101110111010101110111011100110111000101000111011101110111000001000001011001110111001101110111001001000111001100010010011101110111011101110111010100010111011101110010011101110110011100110111011100000100010101110111010101110111001101110001011101110111010001110110011101110111011100010111011101110111011100000010010000100001000101110011011100010111011101100011011101110010011100010001011101110011011101000111011101110111011100000111010101110101",
		"01100111001001110111011100000010001101000101011101110010011101000111011101110111000001110111010101110111011101110001001001110111001101110111011101110111000101110111000101110111011101110101011101110001001001010111010101110111000000000101000001110101011000000000011101110111011101110111000000010111011101110111011100110110011101110101001001100111011101110010011100110100011101110111011001100111011101010111011100100110011101110111001001110111011101110111011101110111000000010010001101110111001001100111011100000000",
		"01000111011101000111011100110000011101000001010000010001011101100111001001110110011101110111001101010110011101000001000001110010010001110111011101110111011101110100000100000111011101110110011101110011011101110111011100110111011101110101000001110111000001110111001001110111011101110001010001110011001101110111001101110001001101110111011101010111011101110101011001110011000001110100010001110111011101110111001001110111011101110111011001010010000101110000001001110111011101110101011101110001011101010111001001110111",
		"01110111011100010000011101110111001000100100001001110010011101110010011001110101011101110111001000000111011101110111010101110111011001110000000001110111010100000111011101110111011101100111011101010111010101110110001101110010011100100111011101010101010101110100001001110111000100110111001001110111011101110111000000100001011101110010011101110111000000010111011101110111000100010000001000110010010101100111001101110111011101110010011101000010000101110111011101110111000101110111011101110111011101110010011101110100",
		"01100111010001110011010101110001011101110101001001110111000001110111011101100100011101110101011101110111011101110111011101110111011100000000000001110000010001010011011101110111000101010100001101010111011001110111010001110111011101110001000100110001011101110010011100100111011100010111011101110111010100000111000101110101000001110111011001100101001101110111011101110111000001110100011101100100011100110111010101110111010101110111001001110111000101110111011101110101001001000111010101110111011101110111011100110111",
		"01110111011101110111000001010000011101110110011101010011011100010111011001110111011101110111011101110111011101110111001001110100001100010111000101010111011001110110001101110000000100100111011100110111011101110111011101010101010000110000011001010111011101110111011101110111011101110110011101110111011101110001011001110100000001100100011101110100000100110001001101110111011101110111011100010111010101100111011101110111011101110010011100010111011101010111011101110001011100110001011101000111011100100111011101110001",
		"01110000000100000111011101110010000101110101010100110111001000000111010001110111011101110111011100000101000001110111011101110100011101110111011101010010011101000011011101110010001101110011011101110011011001110001010001110111011101010111010000100111010001110111011101110111010001110111000100100110011001110000001000100111011101110111011101110010001000000001001001110011011101110111000001110001001101110111011101110111001000110011001001110001000101110100011100000010011101110111010101110011011101110100011100010000",
		"01110111011101110111011100010111011101110011010101000111001100100111001101110111011101000111011101110101000100010111011101110111011101010000000001000000000001100111011101100111011101110111001000000111001001110010010000000111001000110111011101110010011101110010011100110111011101110111000101110111011100010111000001110111011101110111001101110100011001110101011001110111011101110111000101010110011101110001011101110011000100110111010101110111011101110001011101110111011101110001000101110111001001110100011101110111",
		"01010111011100110010011100110111010101100111010100000010000000010111001101010000011101110000011100110111011101000111011101110111010001110101001101110110011101100101011100110111000001110000000101110011001001110001011101000111011101110111011101010111011101110111011101110111001100110100011101110101011101110001000101110111010101110111000101010111011100010011001001110001000101100110011100100000000101110111011100000111011101110111011100000111011101110111011101110110000101100001011100110111001001110111000101000111",
		"01100111011101110001011101010011011100010111010001110111011101110111011101110001001101110111011101110111011101110111011001110111000101110001010001110000011101110001000001110111010001110110011101010110010000010111011101110101011101110010001001110100011000110001011101010001011101110111011100100001010100000011011101110111011101110111011101110010000101110001011100100111000101100111000001110110011101110100010101000101011100010111011101110010011101110110000001110111010101110111011001110111010100110111001001110111",
		"00010111011001010111011100000001011100100010011101110111011101000110000101010100000101110111011001010110010000000111011000110111001001110000000100000111001001110111001001010111010001010101001101000111011101010111011100010111011101110111011101110101001101110111011101110111011101100111011101010110011101110001011101110001011100000111011100010111010000100101011101110010000100010111011101010111011101110111011100010111011101110111011101110101011101110111011101110110010001110011011101110111010101110111011101010000",
		"01010111011101000000000101110001000001110101011100110011001000010111011101010111011100000111011101010001000001000111011101110111011100010111000101110111011100000010000000100111011000100111001101100111001101110011010001100111011101000000011101110111010101010101011100010111001001100111000000110111011101100110011101110100010001110101011101010000011101110111010001010010000101110110011101110010011101110111011101110000000101110111011101000111010101110010011101000000010000100111011101010111010100110111011101110111",
		"01010111001101110111010100100111011101110111011101010111000101110111011001110111011100010111011100000001001001110111001001110111010001110111011101110010011101110000011100110000011101010110001001110111011101110101011100000111011101000100011101110111010000010111011100100011010100110000001000110000011101100010011101110000011101110100011101110100001100110111011100010111011101110000001001110111011101000111001001110111011101110111011101110010011000110111011100110010011100010111010101100111011000100000000100110111",
		"00000000000100110110000101110111011101110000011101110111001101110111010000000001011100000000011101100111011101000111011100110000000000100111011101110111011100000101000001110111011101110111011101110111011101110111011101110111001001010100000001110000011101110111011101110111011101000111011101110111000000000010000101110110001101110001010001110110000000100001001101110100011000010111011101110111011100000111011001010010011100000111001101110001010101110101011100000111000001110111011101000111011101110100011101110111",
		"01110010001101110111011101110111011101110111000000010111011101110010000000000111011101110100010101000000011101000000011101110111011101110101011001010111011001110011011101110111011101110110011101100011011101110111011101110101000100000111011101110111011101110110000101110000000001110111011101110101011100110100001001010111011101110111011101000001011101110010001001110110000001110110011101000111011100110111011101110011011100110100011101110111011101100111001101110111011100100111011101110111001001100101011101110111",
		"01110111011001110111011101110000000001110011011101110111010100100111001001010111011100110011001100010111011101110111011101110100001100000101000000010100011101000001011001110001000000010111011000000100001000000100011101110000011100100111011101010111010001110111011101100010011101110111011100000111010001110111010101000111010101110111011101110001000100110110011101100111011001100111010001110101000101110100011101010000001101100011011101110111010001110001010001010001001001100001011101110111010001110010011001110011",
		"01010111011101110111010100100111011101110111011100010010011101110000011101110001011100000111011100010111011100000111011101110001010101100110011101110111001001110011011101100100011100010111011101110111000101110111011101000111011101110111011100000111011100000000011101000111011001000111011101110101010101110111011101110111010101110111010000100111011101110111011101110111010101110101010101110001000101100111011101110111011101110111011101010111011101110111010101110111011100010111000101110111011101110111011101100110",
		"01110111011101110110011100110111011101110111001100100110011101110111011101110000001001110111011101010111011101110111000001010111011001110011011101110111011101110101011100110001011101110010011101110111011101110111011101110000011101110001000101110110011101110111011101100111001100010111001001110001001101110011011101110010000100110010011100110000011101110010011101110111011100010011011100100111011101110111011101110111001100100111000001110111011101110111011101010001011101000111010101100111010100000111011101010111",
		"01010111010000000000011101110111010000110001011101010111011101110111010000110010011101110000011101110111000000100101011101000111011101100001011101100111011101110111011101110111011101010111011101110111011100010111011101110011011001010111011101110111011101010110011101110111011101100111011001010111001101100101011101110111011001110100011101100111011100000100011100010011001001110111011101110111001001010111001001110111011101110111011101110111000001110111011101010101000001110111001000000111011100110111011101100111",
		"00000111011101110001010001110100011101100111010001110011011101000010000001110011000101110111011101110011011101110101011100010111011101110111011101110111011100100111011101100111011101110111011000100111010101110010011101110111011101110111011100000110011101110011011101110111001101110111001101110111010101110101010101100000011100010111011101110111001101110111011100000000011100100101001001110111011101110110011101110111011101110011010100110110011101100111000101110010011101110111011101010110000001110111011101110111",
		"00110111001101110111011001010101001001110111010101110110011101110111001100100011000001110110011101110111001001110000000101100110011101110111001101100111011101000111011101110111000000100111011100100111011101110111011101110111011101110100010001110110010001110101001101110111011001110111000101110001011101110111011000010101011101110111011101110101011101110110011101010111011001110101011001000011011101110111011101000000000100100111001101110100011101110111001000100111000000100111001101110100011101000000011101110011",
		"01110101011101110111010101100111011001110111010001110111011101110111010001110010011101000110011101010000011101110101001101100111011100110111011000000111011001110111011101110111011101110111010100010111001101000111011101000111000001000111000100010101011100100111001100000111011101110000011001110111011001110111011101110111011100110111001101110011011101110001011101100111011001110111010101110111011100100111011101110111011101000111011100000111001000000001000001100111010101110101001000110111011100100111011101110001",
		"01010111000001000111011100010010010001110111011101110101001101110111001001110000011101110000010101110111011101010110011100110011011101100111011101110111011101110111000100010111001000110010011101000001010101110111011101110111010101110111000001110111011101110011011101110111011101110111010101110111011101110111011100110101011101110111001101110010011101110111011101000111001000110111011101110001001101110111011101110111011101110000010101110011010000100111011101110111010101110111010001110000000100000111001100000111",
		"01110101011000100100001101110001011101110111011101000111011101110010010001110011001100010101010001010111011101110111000000000111010100000111001001000111010001110111011100010000010000100010011101010111010101110111011100000010011101110000011101110111011101110110011101110011011001110111010001110111000000110010011101110111011101110100010101110111000101110111011101110111011101110111010001110101011101110111011101010111011100100111011101110111011101110001011101110111011101110111011101110111010001110101011001110100",
		"00100111011100010011011101110111011100010001000100110111011101110111011101110111000101110011011101110111011100010111001101110110011100100001011101110011010100100101011101110100001100100010010101010111011100010111011100110000011101110111011100000110010001110110011101110111011101110110001001110101011000010111011100110111001001110111011101110101000001000111011100010111011000110100011101110111001101110111011100000101011101110001000100010111011101110111011101110101011101110011000101110111011101110111011101110111",
		"01110101011101000111001101100011011100100011010001110000001101110111010001110001011100100000011101110111011101010001001101110110010101110111000001110010011101110111011101110101011101110111001101110000011101110110001001000111011101110011000101110111001101110111000001100010011100100111011101000111011101110111011101110110011001110111011101010111010100100000001101110111011101010111011101110111010100100111011101110111011100000111011101110001000101110010011100010100011101110111011101110000011101110111000001000000",
		"01100111011101110111011100110111001001110111011100010011001101110010011101110100001101110010011101110000011101010111011101000111000001010001010101010111011101010111011101110111011100000111011101110111010001110111010101010111011100100011011000110111001001000111011101110110011101110011011001110111011101110111011100110100011001110101010100000100010001110111011001110111000001110111011101010101011100110111011101110111011100010011001101110111011000100111001001110011011101110010010001110101011101110001011101110111",
		"01110111011101000111011101110111011101010111010001110001011101110111011101110111011101110000011100010111011101110110010100100110001000010000011101110000001101000110000001010011011101110111011101110110001001010010011101000111011101110111011100010111011101110111011101000111011100100111011101000010000001100011001000100111000001100111011101110000011101110010010001000111011101110111011001110111000001110111010000010111011101110111011100110110000100000111011101110001011101110111001101110111011101110111010101110111",
		"00110001011100000111011100000111011100010101001001110111011101110111011101110010011101110111010100110010011101110110001101110111011101110111011101010000010000110000001001110111000101000000011101110111011101100111011101110000011101100111010001110111011100110100010001110111001101010111011100100100010101110100011100000111010001110111000001110111011101110111011101110111011101000110011000000111011101100101011100010011010000110010011001110100011101110011011101110001011101110100011101110110001101100110001100000110",
		"01110111011101110010011100010111000101100111011100100111011101110111011101110111000100010001001101110001010000100111000101110111011101110011011101100101011101010111001001110111011101110100010101110000011101100000011100110111011100000111011101110110011101110011011101110001001100000111011101110111011101110111010001110111001001110111011101010111011001100111000001110111011101110110001000010111011101000111011101110111011101110000011100110111001001000000010001110101011100110111011100110010011101110111011101010001",
		"00110111011101110111000000000111011101110101011101010011011100010001000001000111011101110100011101000001011001100111011101110111011101000011001100110111010100000000011001100111011101100001000101100111011101100111010101110111001001110101001101100111001101110111011101110111011101100111010001110111000001110111011101110111000001110111011101010101011101110110011101110011011101100111011101110100011100000010011101110100011101010111000001000011011100010111011101110000011100100001011101110111011100010111011101110101",
		"00100010011101110001000101110110011101000001011101110111011100110001000001000101011101110111011101010011011100000111011101110000011100110111000000010111011101110001011101110000011101110111001001110010000001110010011101110000000101110111011101010101011101110111001000010111000001110111000001110111011101110111011101110111011100010111011101110110001101110111011101000100011101110101011101110111011101110001011101110000011101110101000101110010010001100101011101110111011101110101011101110111011001000010011100010001",
		"00110010011100010000010001110111010000000111001000000010011001100111010001110110000101110000001000100111010001110011011001110100011100110110011101110111011101110111011101000111011101000010011100110111011101110010011100100100001100100111011101010111011101110111011100110001011001110011011100010111011101110100011100000111011101110111001001110100010001110011011101000000011101110111001101110011001101110001010100100100011001110101011100110111011101110111011101110111011101110100001001110111000000010001010000000000"
	);

begin

	rom_behavior	: process(clka)
	begin

		if clka'event and clka = '1'
		then

			douta <= mem(to_integer(unsigned(addra)));

		end if;

	end process rom_behavior;

end architecture behavior;

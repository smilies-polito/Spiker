library ieee;
use ieee.std_logic_1164.all;


entity lfsr is

end entity lfsr;


architecture behaviour of lfsr is

begin

end architecture behaviour;

library ieee;
use ieee.std_logic_1164.all;


--  RAMB36E1   : In order to incorporate this function into the design,
--    VHDL     : the following instance declaration needs to be placed
--  instance   : in the body of the design code.  The instance name
-- declaration : (RAMB36E1_inst) and/or the port declarations after the
--    code     : "=>" declaration maybe changed to properly reference and
--             : connect this function to the design.  All inputs and outputs
--             : must be connected.

--   Library   : In addition to adding the instance declaration, a use
-- declaration : statement for the UNISIM.vcomponents library needs to be
--     for     : added before the entity declaration.  This library
--   Xilinx    : contains the component declarations for all Xilinx
-- primitives  : primitives and points to the models that will be used
--             : for simulation.

--  Copy the following two statements and paste them before the
--  Entity declaration, unless they already exist.

library UNISIM;
use UNISIM.vcomponents.all;


entity bram_sdp is

	port(
		-- input
		clk		: in std_logic;
		di		: in std_logic_vector(71 downto 0);
		rdaddr		: in std_logic_vector(15 downto 0);
		rden		: in std_logic;
		wraddr		: in std_logic_vector(15 downto 0);
		wren		: in std_logic;

		-- output
		do		: out std_logic_vector(71 downto 0)
				
	);

end entity bram_sdp;


architecture behaviour of bram_sdp is

begin


	-- RAMB36E1: 36K-bit Configurable Synchronous Block RAM
	--           Artix-7
	-- Xilinx HDL Language Template, version 2020.2

	RAMB36E1_inst : RAMB36E1
		generic map (
			-- Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
			RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
			-- Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
			SIM_COLLISION_CHECK => "ALL",
			-- DOA_REG, DOB_REG: Optional output register (0 or 1)
			DOA_REG => 0,
			DOB_REG => 0,
			EN_ECC_READ => FALSE,                                                            -- Enable ECC decoder,
												       -- FALSE, TRUE
			EN_ECC_WRITE => FALSE,                                                           -- Enable ECC encoder,
												       -- FALSE, TRUE
			-- INITP_00 to INITP_0F: Initial contents of the parity memory array
			INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			-- INIT_00 to INIT_7F: Initial contents of the data memory array
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
			-- INIT_A, INIT_B: Initial values on output ports
			INIT_A => X"000000000",
			INIT_B => X"000000000",
			-- Initialization File: RAM initialization file
			INIT_FILE => "NONE",
			-- RAM Mode: "SDP" or "TDP" 
			RAM_MODE => "SDP",
			-- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
			RAM_EXTENSION_A => "NONE",
			RAM_EXTENSION_B => "NONE",
			-- READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
			READ_WIDTH_A => 0,                                                               -- 0-72
			READ_WIDTH_B => 0,                                                               -- 0-36
			WRITE_WIDTH_A => 0,                                                              -- 0-36
			WRITE_WIDTH_B => 0,                                                              -- 0-72
			-- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
			RSTREG_PRIORITY_A => "RSTREG",
			RSTREG_PRIORITY_B => "RSTREG",
			-- SRVAL_A, SRVAL_B: Set/reset value for output
			SRVAL_A => X"000000000",
			SRVAL_B => X"000000000",
			-- Simulation Device: Must be set to "7SERIES" for simulation behavior
			SIM_DEVICE => "7SERIES",
			-- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
			WRITE_MODE_A => "WRITE_FIRST",
			WRITE_MODE_B => "WRITE_FIRST" 
		)

		port map (
			-- Cascade Signals: 1-bit (each) output: BRAM cascade ports (to create 64kx1)
			CASCADEOUTA => open,     -- 1-bit output: A port cascade
			CASCADEOUTB => open,     -- 1-bit output: B port cascade
			-- ECC Signals: 1-bit (each) output: Error Correction Circuitry ports
			DBITERR => open,             -- 1-bit output: Double bit error status
			ECCPARITY => open,         -- 8-bit output: Generated error correction parity
			RDADDRECC => open,         -- 9-bit output: ECC read address
			SBITERR => open,             -- 1-bit output: Single bit error status
			-- Port A Data: 32-bit (each) output: Port A data
			DOADO => do(39 downto 8),                 -- 32-bit output: A port data/LSB data
			DOPADOP => do(3 downto 0),             -- 4-bit output: A port parity/LSB parity
			-- Port B Data: 32-bit (each) output: Port B data
			DOBDO => do(71 downto 40),                 -- 32-bit output: B port data/MSB data
			DOPBDOP => do(7 downto 4),             -- 4-bit output: B port parity/MSB parity
			-- Cascade Signals: 1-bit (each) input: BRAM cascade ports (to create 64kx1)
			CASCADEINA => '0',       -- 1-bit input: A port cascade
			CASCADEINB => '0',       -- 1-bit input: B port cascade
			-- ECC Signals: 1-bit (each) input: Error Correction Circuitry ports
			INJECTDBITERR => '0', -- 1-bit input: Inject a double bit error
			INJECTSBITERR => '0', -- 1-bit input: Inject a single bit error

			-- Port A Address/Control Signals: 16-bit (each) input: Port A address and control signals (read port
			-- when RAM_MODE="SDP")
			ADDRARDADDR => rdaddr,     -- 16-bit input: A port address/Read address
			CLKARDCLK => clk,         -- 1-bit input: A port clock/Read clock
			ENARDEN => rden,             -- 1-bit input: A port enable/Read enable
			REGCEAREGCE => '0',     -- 1-bit input: A port register enable/Register enable
			RSTRAMARSTRAM => '0', -- 1-bit input: A port set/reset
			RSTREGARSTREG => '0', -- 1-bit input: A port register set/reset
			WEA => (others => '0'),                     -- 4-bit input: A port write enable

			-- Port A Data: 32-bit (each) input: Port A data
			DIADI => di(39 downto 8),                 -- 32-bit input: A port data/LSB data
			DIPADIP => di(3 downto 0),             -- 4-bit input: A port parity/LSB parity
			-- Port B Address/Control Signals: 16-bit (each) input: Port B address and control signals (write port
			-- when RAM_MODE="SDP")
			ADDRBWRADDR => wraddr,     -- 16-bit input: B port address/Write address
			CLKBWRCLK => clk,         -- 1-bit input: B port clock/Write clock
			ENBWREN => wren,             -- 1-bit input: B port enable/Write enable
			REGCEB => '0',               -- 1-bit input: B port register enable
			RSTRAMB => '0',             -- 1-bit input: B port set/reset
			RSTREGB => '0',             -- 1-bit input: B port register set/reset
			WEBWE => (others => '0'),                 -- 8-bit input: B port write enable/Write enable
			-- Port B Data: 32-bit (each) input: Port B data
			DIBDI => di(71 downto 40),                 -- 32-bit input: B port data/MSB data
			DIPBDIP => di(7 downto 4)              -- 4-bit input: B port parity/MSB parity
		);

					
end architecture behaviour;	

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_128x10_exc_ip is
	port(
		clka	: in std_logic;
		addra	: in std_logic_vector(6 downto 0);
		douta	: out std_logic_vector(39 downto 0)
	);
end entity rom_128x10_exc_ip; 

architecture behavior of rom_128x10_exc_ip is

	type rom_type is array(0 to 127) of std_logic_vector(39 downto 0);

	constant mem	: rom_type := (
		"0111000101110101001001110011010001110111",
		"0111001001110101011101000100011101110111",
		"0111011101110000011101010011011101110111",
		"0000000101110111001100100111001001010111",
		"0011011100000111011101100101001000010111",
		"0001011001110111000000010011001100110111",
		"0101000001000011000001110111011101110111",
		"0001000001110001011001110011011101110111",
		"0000011101110011000000000110011101110111",
		"0101011100110001000001010111010001110100",
		"0100011101110010011001010111011101110111",
		"0010011101110111001101110100010101110111",
		"0111011101010111011101110111011101110111",
		"0000011101110111011100100111011100110011",
		"0000010101110011011101110111011001000101",
		"0011011000000111011001110111011101110111",
		"0011011101110111011101110011011100110101",
		"0000011101110101011101110111011101110001",
		"0101000101110000000101000011011101110111",
		"0101011101110100011101110111011101110001",
		"0011011100000100000001110111001000110111",
		"0101011101110110011101110000001001010010",
		"0001011101110111011101110101011101110111",
		"0011011101100111001101110011001001010010",
		"0010011101110111000101000110010100010111",
		"0111000001110111011100010111010100110111",
		"0101010101110110011101110101011100000110",
		"0111010101110001011101000101011100110010",
		"0111000100000011011101000010011101110010",
		"0100011101110101011100110111011101110111",
		"0111001001110111011101110111011101110101",
		"0111011101000111011101110111011101110111",
		"0111010101110111010000000111001101010111",
		"0111010101110011011101110111001101110110",
		"0111011101110111011101010010011101000111",
		"0111011100010111011101110101010001110111",
		"0111001001110110011001100111010101000111",
		"0111001100100111011100110011010101000111",
		"0111010001010111000100110000011100100010",
		"0111011100110111011101010100011101110000",
		"0101010001110111011101110111011101010101",
		"0111001101100111011101110111010100110110",
		"0111011101110111011001110100000001000111",
		"0010011101110111011101110001010000010100",
		"0111000001110111011101010110010001000111",
		"0111011100000111011101010111011101010111",
		"0111010101110010001101110011011101100111",
		"0111011101110111000000110111011100100001",
		"0111000001110101011101110111011101110101",
		"0111011000110101000001010111011101000100",
		"0111011101110011011101110011011101110111",
		"0110011101110101001100110001011100010111",
		"0010011101110001011101110111011101110100",
		"0011010101110110010001110000001101110111",
		"0000011101000001011101110010011101000111",
		"0111011101110111011101110111011101110010",
		"0010000101100111000001110111011101110001",
		"0100011000010111000101110111010001110111",
		"0111010101110111011100100111010101110111",
		"0100011100010101011101010111000000010110",
		"0111011101100111011101110111000001110110",
		"0010011101110111011100000010000001110001",
		"0011000101100111011101110110010101010010",
		"0110011101110111000001110010011101110011",
		"0111011101110101001101110111011101110111",
		"0111000001110111010000010111011101110111",
		"0010011100110111011100100111010101110011",
		"0110011100100111010001110011011101110111",
		"0111010100100111011101110111011100000111",
		"0010000100010111001001110111010001010111",
		"0111011101110111010001110000000100100111",
		"0111011001110011000101000111011101110010",
		"0111011100010111001101110111000100010111",
		"0111000100100111000101000101011101110011",
		"0111011101110111011101110010000100000111",
		"0001011101110111011101110111010000000111",
		"0111000101000000011101110011011101000111",
		"0111010001110001010101110111010100010110",
		"0110011101110111010001110000010101110111",
		"0111011101110001011101110010011101110011",
		"0111000001110001011101110111010000100111",
		"0101011001110100000001110111000001110000",
		"0001010001100111011101110111000000000010",
		"0111011101110111011101110111011001110111",
		"0100010101110111011101110111011101110000",
		"0111011101110100011100100101010101000011",
		"0011011101000111010001110101011101100011",
		"0111001001110000011101010111011101110011",
		"0100011101100111011101010000011000100111",
		"0001010000110111011101000111010001110111",
		"0000011101110111000101000000011101110001",
		"0111000001100110000001010000000001110101",
		"0111011101110011001000000111010000000111",
		"0111001101110001011001110111010101110111",
		"0011001001110111011100000001001001110100",
		"0111011101110100001001110111011101110100",
		"0111010101110111011101010001011101100111",
		"0000011101100111011101110100011101110111",
		"0000011101110011011101110111011101110111",
		"0111011101010111011101110100011000010111",
		"0111011001010111011101000011011101110111",
		"0111011101110111011101010110011101110011",
		"0110011101110011011100110111001001100101",
		"0111011101110111011101110001011101110111",
		"0010010001110111011101110111011100000011",
		"0111011001110111011001010111011101100111",
		"0111011100110111011101110101010101110111",
		"0000011100110111011001110111011101110111",
		"0111011101110111010001110111011101110111",
		"0000000000100000011101100000011101110110",
		"0001011101110111011101110111011101110010",
		"0110011101110101011001110111000001100111",
		"0110000100100111011101000000011001110111",
		"0101011101110111010000110111011100110001",
		"0111011101110010011100100111000101110111",
		"0011011101000111011101110010011101110000",
		"0000011000110111001001110000011100100111",
		"0011001101110111011100110101011101110110",
		"0111000001110111011001110100011100000010",
		"0110011001000010011101000001011101110111",
		"0001011101110111000101000001011101110011",
		"0111011101110011011101110111011101110111",
		"0111011001110111010001110111011101010111",
		"0111011101110111011101110000010001000111",
		"0111001101110111011100100111010101000001",
		"0111011101110111011100000010000001110110",
		"0111000001110111010001010111010000000111",
		"0110000000010011001001110110000100000111"
	);

begin

	rom_behavior	: process(clka)
	begin

		if clka'event and clka = '1'
		then

			douta <= mem(to_integer(unsigned(addra)));

		end if;

	end process rom_behavior;

end architecture behavior;

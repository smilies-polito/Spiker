library ieee;
use ieee.std_logic_1164.all;

entity input_interface is

end entity input_interface;

architecture behaviour of input_interface is
begin

end architecture behaviour;

---------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or
-- distribute this software, either in source code form or as a compiled
-- binary, for any purpose, commercial or non-commercial, and by any
-- means.
--
-- In jurisdictions that recognize copyright laws, the author or authors
-- of this software dedicate any and all copyright interest in the
-- software to the public domain. We make this dedication for the benefit
-- of the public at large and to the detriment of our heirs and
-- successors. We intend this dedication to be an overt act of
-- relinquishment in perpetuity of all present and future rights to this
-- software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR
-- OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE.
--
-- For more information, please refer to <http://unlicense.org/>
---------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;


entity mux_1024to1 is
    port (
        mux_sel : in std_logic_vector(9 downto 0);
        in0 : in std_logic;
        in1 : in std_logic;
        in2 : in std_logic;
        in3 : in std_logic;
        in4 : in std_logic;
        in5 : in std_logic;
        in6 : in std_logic;
        in7 : in std_logic;
        in8 : in std_logic;
        in9 : in std_logic;
        in10 : in std_logic;
        in11 : in std_logic;
        in12 : in std_logic;
        in13 : in std_logic;
        in14 : in std_logic;
        in15 : in std_logic;
        in16 : in std_logic;
        in17 : in std_logic;
        in18 : in std_logic;
        in19 : in std_logic;
        in20 : in std_logic;
        in21 : in std_logic;
        in22 : in std_logic;
        in23 : in std_logic;
        in24 : in std_logic;
        in25 : in std_logic;
        in26 : in std_logic;
        in27 : in std_logic;
        in28 : in std_logic;
        in29 : in std_logic;
        in30 : in std_logic;
        in31 : in std_logic;
        in32 : in std_logic;
        in33 : in std_logic;
        in34 : in std_logic;
        in35 : in std_logic;
        in36 : in std_logic;
        in37 : in std_logic;
        in38 : in std_logic;
        in39 : in std_logic;
        in40 : in std_logic;
        in41 : in std_logic;
        in42 : in std_logic;
        in43 : in std_logic;
        in44 : in std_logic;
        in45 : in std_logic;
        in46 : in std_logic;
        in47 : in std_logic;
        in48 : in std_logic;
        in49 : in std_logic;
        in50 : in std_logic;
        in51 : in std_logic;
        in52 : in std_logic;
        in53 : in std_logic;
        in54 : in std_logic;
        in55 : in std_logic;
        in56 : in std_logic;
        in57 : in std_logic;
        in58 : in std_logic;
        in59 : in std_logic;
        in60 : in std_logic;
        in61 : in std_logic;
        in62 : in std_logic;
        in63 : in std_logic;
        in64 : in std_logic;
        in65 : in std_logic;
        in66 : in std_logic;
        in67 : in std_logic;
        in68 : in std_logic;
        in69 : in std_logic;
        in70 : in std_logic;
        in71 : in std_logic;
        in72 : in std_logic;
        in73 : in std_logic;
        in74 : in std_logic;
        in75 : in std_logic;
        in76 : in std_logic;
        in77 : in std_logic;
        in78 : in std_logic;
        in79 : in std_logic;
        in80 : in std_logic;
        in81 : in std_logic;
        in82 : in std_logic;
        in83 : in std_logic;
        in84 : in std_logic;
        in85 : in std_logic;
        in86 : in std_logic;
        in87 : in std_logic;
        in88 : in std_logic;
        in89 : in std_logic;
        in90 : in std_logic;
        in91 : in std_logic;
        in92 : in std_logic;
        in93 : in std_logic;
        in94 : in std_logic;
        in95 : in std_logic;
        in96 : in std_logic;
        in97 : in std_logic;
        in98 : in std_logic;
        in99 : in std_logic;
        in100 : in std_logic;
        in101 : in std_logic;
        in102 : in std_logic;
        in103 : in std_logic;
        in104 : in std_logic;
        in105 : in std_logic;
        in106 : in std_logic;
        in107 : in std_logic;
        in108 : in std_logic;
        in109 : in std_logic;
        in110 : in std_logic;
        in111 : in std_logic;
        in112 : in std_logic;
        in113 : in std_logic;
        in114 : in std_logic;
        in115 : in std_logic;
        in116 : in std_logic;
        in117 : in std_logic;
        in118 : in std_logic;
        in119 : in std_logic;
        in120 : in std_logic;
        in121 : in std_logic;
        in122 : in std_logic;
        in123 : in std_logic;
        in124 : in std_logic;
        in125 : in std_logic;
        in126 : in std_logic;
        in127 : in std_logic;
        in128 : in std_logic;
        in129 : in std_logic;
        in130 : in std_logic;
        in131 : in std_logic;
        in132 : in std_logic;
        in133 : in std_logic;
        in134 : in std_logic;
        in135 : in std_logic;
        in136 : in std_logic;
        in137 : in std_logic;
        in138 : in std_logic;
        in139 : in std_logic;
        in140 : in std_logic;
        in141 : in std_logic;
        in142 : in std_logic;
        in143 : in std_logic;
        in144 : in std_logic;
        in145 : in std_logic;
        in146 : in std_logic;
        in147 : in std_logic;
        in148 : in std_logic;
        in149 : in std_logic;
        in150 : in std_logic;
        in151 : in std_logic;
        in152 : in std_logic;
        in153 : in std_logic;
        in154 : in std_logic;
        in155 : in std_logic;
        in156 : in std_logic;
        in157 : in std_logic;
        in158 : in std_logic;
        in159 : in std_logic;
        in160 : in std_logic;
        in161 : in std_logic;
        in162 : in std_logic;
        in163 : in std_logic;
        in164 : in std_logic;
        in165 : in std_logic;
        in166 : in std_logic;
        in167 : in std_logic;
        in168 : in std_logic;
        in169 : in std_logic;
        in170 : in std_logic;
        in171 : in std_logic;
        in172 : in std_logic;
        in173 : in std_logic;
        in174 : in std_logic;
        in175 : in std_logic;
        in176 : in std_logic;
        in177 : in std_logic;
        in178 : in std_logic;
        in179 : in std_logic;
        in180 : in std_logic;
        in181 : in std_logic;
        in182 : in std_logic;
        in183 : in std_logic;
        in184 : in std_logic;
        in185 : in std_logic;
        in186 : in std_logic;
        in187 : in std_logic;
        in188 : in std_logic;
        in189 : in std_logic;
        in190 : in std_logic;
        in191 : in std_logic;
        in192 : in std_logic;
        in193 : in std_logic;
        in194 : in std_logic;
        in195 : in std_logic;
        in196 : in std_logic;
        in197 : in std_logic;
        in198 : in std_logic;
        in199 : in std_logic;
        in200 : in std_logic;
        in201 : in std_logic;
        in202 : in std_logic;
        in203 : in std_logic;
        in204 : in std_logic;
        in205 : in std_logic;
        in206 : in std_logic;
        in207 : in std_logic;
        in208 : in std_logic;
        in209 : in std_logic;
        in210 : in std_logic;
        in211 : in std_logic;
        in212 : in std_logic;
        in213 : in std_logic;
        in214 : in std_logic;
        in215 : in std_logic;
        in216 : in std_logic;
        in217 : in std_logic;
        in218 : in std_logic;
        in219 : in std_logic;
        in220 : in std_logic;
        in221 : in std_logic;
        in222 : in std_logic;
        in223 : in std_logic;
        in224 : in std_logic;
        in225 : in std_logic;
        in226 : in std_logic;
        in227 : in std_logic;
        in228 : in std_logic;
        in229 : in std_logic;
        in230 : in std_logic;
        in231 : in std_logic;
        in232 : in std_logic;
        in233 : in std_logic;
        in234 : in std_logic;
        in235 : in std_logic;
        in236 : in std_logic;
        in237 : in std_logic;
        in238 : in std_logic;
        in239 : in std_logic;
        in240 : in std_logic;
        in241 : in std_logic;
        in242 : in std_logic;
        in243 : in std_logic;
        in244 : in std_logic;
        in245 : in std_logic;
        in246 : in std_logic;
        in247 : in std_logic;
        in248 : in std_logic;
        in249 : in std_logic;
        in250 : in std_logic;
        in251 : in std_logic;
        in252 : in std_logic;
        in253 : in std_logic;
        in254 : in std_logic;
        in255 : in std_logic;
        in256 : in std_logic;
        in257 : in std_logic;
        in258 : in std_logic;
        in259 : in std_logic;
        in260 : in std_logic;
        in261 : in std_logic;
        in262 : in std_logic;
        in263 : in std_logic;
        in264 : in std_logic;
        in265 : in std_logic;
        in266 : in std_logic;
        in267 : in std_logic;
        in268 : in std_logic;
        in269 : in std_logic;
        in270 : in std_logic;
        in271 : in std_logic;
        in272 : in std_logic;
        in273 : in std_logic;
        in274 : in std_logic;
        in275 : in std_logic;
        in276 : in std_logic;
        in277 : in std_logic;
        in278 : in std_logic;
        in279 : in std_logic;
        in280 : in std_logic;
        in281 : in std_logic;
        in282 : in std_logic;
        in283 : in std_logic;
        in284 : in std_logic;
        in285 : in std_logic;
        in286 : in std_logic;
        in287 : in std_logic;
        in288 : in std_logic;
        in289 : in std_logic;
        in290 : in std_logic;
        in291 : in std_logic;
        in292 : in std_logic;
        in293 : in std_logic;
        in294 : in std_logic;
        in295 : in std_logic;
        in296 : in std_logic;
        in297 : in std_logic;
        in298 : in std_logic;
        in299 : in std_logic;
        in300 : in std_logic;
        in301 : in std_logic;
        in302 : in std_logic;
        in303 : in std_logic;
        in304 : in std_logic;
        in305 : in std_logic;
        in306 : in std_logic;
        in307 : in std_logic;
        in308 : in std_logic;
        in309 : in std_logic;
        in310 : in std_logic;
        in311 : in std_logic;
        in312 : in std_logic;
        in313 : in std_logic;
        in314 : in std_logic;
        in315 : in std_logic;
        in316 : in std_logic;
        in317 : in std_logic;
        in318 : in std_logic;
        in319 : in std_logic;
        in320 : in std_logic;
        in321 : in std_logic;
        in322 : in std_logic;
        in323 : in std_logic;
        in324 : in std_logic;
        in325 : in std_logic;
        in326 : in std_logic;
        in327 : in std_logic;
        in328 : in std_logic;
        in329 : in std_logic;
        in330 : in std_logic;
        in331 : in std_logic;
        in332 : in std_logic;
        in333 : in std_logic;
        in334 : in std_logic;
        in335 : in std_logic;
        in336 : in std_logic;
        in337 : in std_logic;
        in338 : in std_logic;
        in339 : in std_logic;
        in340 : in std_logic;
        in341 : in std_logic;
        in342 : in std_logic;
        in343 : in std_logic;
        in344 : in std_logic;
        in345 : in std_logic;
        in346 : in std_logic;
        in347 : in std_logic;
        in348 : in std_logic;
        in349 : in std_logic;
        in350 : in std_logic;
        in351 : in std_logic;
        in352 : in std_logic;
        in353 : in std_logic;
        in354 : in std_logic;
        in355 : in std_logic;
        in356 : in std_logic;
        in357 : in std_logic;
        in358 : in std_logic;
        in359 : in std_logic;
        in360 : in std_logic;
        in361 : in std_logic;
        in362 : in std_logic;
        in363 : in std_logic;
        in364 : in std_logic;
        in365 : in std_logic;
        in366 : in std_logic;
        in367 : in std_logic;
        in368 : in std_logic;
        in369 : in std_logic;
        in370 : in std_logic;
        in371 : in std_logic;
        in372 : in std_logic;
        in373 : in std_logic;
        in374 : in std_logic;
        in375 : in std_logic;
        in376 : in std_logic;
        in377 : in std_logic;
        in378 : in std_logic;
        in379 : in std_logic;
        in380 : in std_logic;
        in381 : in std_logic;
        in382 : in std_logic;
        in383 : in std_logic;
        in384 : in std_logic;
        in385 : in std_logic;
        in386 : in std_logic;
        in387 : in std_logic;
        in388 : in std_logic;
        in389 : in std_logic;
        in390 : in std_logic;
        in391 : in std_logic;
        in392 : in std_logic;
        in393 : in std_logic;
        in394 : in std_logic;
        in395 : in std_logic;
        in396 : in std_logic;
        in397 : in std_logic;
        in398 : in std_logic;
        in399 : in std_logic;
        in400 : in std_logic;
        in401 : in std_logic;
        in402 : in std_logic;
        in403 : in std_logic;
        in404 : in std_logic;
        in405 : in std_logic;
        in406 : in std_logic;
        in407 : in std_logic;
        in408 : in std_logic;
        in409 : in std_logic;
        in410 : in std_logic;
        in411 : in std_logic;
        in412 : in std_logic;
        in413 : in std_logic;
        in414 : in std_logic;
        in415 : in std_logic;
        in416 : in std_logic;
        in417 : in std_logic;
        in418 : in std_logic;
        in419 : in std_logic;
        in420 : in std_logic;
        in421 : in std_logic;
        in422 : in std_logic;
        in423 : in std_logic;
        in424 : in std_logic;
        in425 : in std_logic;
        in426 : in std_logic;
        in427 : in std_logic;
        in428 : in std_logic;
        in429 : in std_logic;
        in430 : in std_logic;
        in431 : in std_logic;
        in432 : in std_logic;
        in433 : in std_logic;
        in434 : in std_logic;
        in435 : in std_logic;
        in436 : in std_logic;
        in437 : in std_logic;
        in438 : in std_logic;
        in439 : in std_logic;
        in440 : in std_logic;
        in441 : in std_logic;
        in442 : in std_logic;
        in443 : in std_logic;
        in444 : in std_logic;
        in445 : in std_logic;
        in446 : in std_logic;
        in447 : in std_logic;
        in448 : in std_logic;
        in449 : in std_logic;
        in450 : in std_logic;
        in451 : in std_logic;
        in452 : in std_logic;
        in453 : in std_logic;
        in454 : in std_logic;
        in455 : in std_logic;
        in456 : in std_logic;
        in457 : in std_logic;
        in458 : in std_logic;
        in459 : in std_logic;
        in460 : in std_logic;
        in461 : in std_logic;
        in462 : in std_logic;
        in463 : in std_logic;
        in464 : in std_logic;
        in465 : in std_logic;
        in466 : in std_logic;
        in467 : in std_logic;
        in468 : in std_logic;
        in469 : in std_logic;
        in470 : in std_logic;
        in471 : in std_logic;
        in472 : in std_logic;
        in473 : in std_logic;
        in474 : in std_logic;
        in475 : in std_logic;
        in476 : in std_logic;
        in477 : in std_logic;
        in478 : in std_logic;
        in479 : in std_logic;
        in480 : in std_logic;
        in481 : in std_logic;
        in482 : in std_logic;
        in483 : in std_logic;
        in484 : in std_logic;
        in485 : in std_logic;
        in486 : in std_logic;
        in487 : in std_logic;
        in488 : in std_logic;
        in489 : in std_logic;
        in490 : in std_logic;
        in491 : in std_logic;
        in492 : in std_logic;
        in493 : in std_logic;
        in494 : in std_logic;
        in495 : in std_logic;
        in496 : in std_logic;
        in497 : in std_logic;
        in498 : in std_logic;
        in499 : in std_logic;
        in500 : in std_logic;
        in501 : in std_logic;
        in502 : in std_logic;
        in503 : in std_logic;
        in504 : in std_logic;
        in505 : in std_logic;
        in506 : in std_logic;
        in507 : in std_logic;
        in508 : in std_logic;
        in509 : in std_logic;
        in510 : in std_logic;
        in511 : in std_logic;
        in512 : in std_logic;
        in513 : in std_logic;
        in514 : in std_logic;
        in515 : in std_logic;
        in516 : in std_logic;
        in517 : in std_logic;
        in518 : in std_logic;
        in519 : in std_logic;
        in520 : in std_logic;
        in521 : in std_logic;
        in522 : in std_logic;
        in523 : in std_logic;
        in524 : in std_logic;
        in525 : in std_logic;
        in526 : in std_logic;
        in527 : in std_logic;
        in528 : in std_logic;
        in529 : in std_logic;
        in530 : in std_logic;
        in531 : in std_logic;
        in532 : in std_logic;
        in533 : in std_logic;
        in534 : in std_logic;
        in535 : in std_logic;
        in536 : in std_logic;
        in537 : in std_logic;
        in538 : in std_logic;
        in539 : in std_logic;
        in540 : in std_logic;
        in541 : in std_logic;
        in542 : in std_logic;
        in543 : in std_logic;
        in544 : in std_logic;
        in545 : in std_logic;
        in546 : in std_logic;
        in547 : in std_logic;
        in548 : in std_logic;
        in549 : in std_logic;
        in550 : in std_logic;
        in551 : in std_logic;
        in552 : in std_logic;
        in553 : in std_logic;
        in554 : in std_logic;
        in555 : in std_logic;
        in556 : in std_logic;
        in557 : in std_logic;
        in558 : in std_logic;
        in559 : in std_logic;
        in560 : in std_logic;
        in561 : in std_logic;
        in562 : in std_logic;
        in563 : in std_logic;
        in564 : in std_logic;
        in565 : in std_logic;
        in566 : in std_logic;
        in567 : in std_logic;
        in568 : in std_logic;
        in569 : in std_logic;
        in570 : in std_logic;
        in571 : in std_logic;
        in572 : in std_logic;
        in573 : in std_logic;
        in574 : in std_logic;
        in575 : in std_logic;
        in576 : in std_logic;
        in577 : in std_logic;
        in578 : in std_logic;
        in579 : in std_logic;
        in580 : in std_logic;
        in581 : in std_logic;
        in582 : in std_logic;
        in583 : in std_logic;
        in584 : in std_logic;
        in585 : in std_logic;
        in586 : in std_logic;
        in587 : in std_logic;
        in588 : in std_logic;
        in589 : in std_logic;
        in590 : in std_logic;
        in591 : in std_logic;
        in592 : in std_logic;
        in593 : in std_logic;
        in594 : in std_logic;
        in595 : in std_logic;
        in596 : in std_logic;
        in597 : in std_logic;
        in598 : in std_logic;
        in599 : in std_logic;
        in600 : in std_logic;
        in601 : in std_logic;
        in602 : in std_logic;
        in603 : in std_logic;
        in604 : in std_logic;
        in605 : in std_logic;
        in606 : in std_logic;
        in607 : in std_logic;
        in608 : in std_logic;
        in609 : in std_logic;
        in610 : in std_logic;
        in611 : in std_logic;
        in612 : in std_logic;
        in613 : in std_logic;
        in614 : in std_logic;
        in615 : in std_logic;
        in616 : in std_logic;
        in617 : in std_logic;
        in618 : in std_logic;
        in619 : in std_logic;
        in620 : in std_logic;
        in621 : in std_logic;
        in622 : in std_logic;
        in623 : in std_logic;
        in624 : in std_logic;
        in625 : in std_logic;
        in626 : in std_logic;
        in627 : in std_logic;
        in628 : in std_logic;
        in629 : in std_logic;
        in630 : in std_logic;
        in631 : in std_logic;
        in632 : in std_logic;
        in633 : in std_logic;
        in634 : in std_logic;
        in635 : in std_logic;
        in636 : in std_logic;
        in637 : in std_logic;
        in638 : in std_logic;
        in639 : in std_logic;
        in640 : in std_logic;
        in641 : in std_logic;
        in642 : in std_logic;
        in643 : in std_logic;
        in644 : in std_logic;
        in645 : in std_logic;
        in646 : in std_logic;
        in647 : in std_logic;
        in648 : in std_logic;
        in649 : in std_logic;
        in650 : in std_logic;
        in651 : in std_logic;
        in652 : in std_logic;
        in653 : in std_logic;
        in654 : in std_logic;
        in655 : in std_logic;
        in656 : in std_logic;
        in657 : in std_logic;
        in658 : in std_logic;
        in659 : in std_logic;
        in660 : in std_logic;
        in661 : in std_logic;
        in662 : in std_logic;
        in663 : in std_logic;
        in664 : in std_logic;
        in665 : in std_logic;
        in666 : in std_logic;
        in667 : in std_logic;
        in668 : in std_logic;
        in669 : in std_logic;
        in670 : in std_logic;
        in671 : in std_logic;
        in672 : in std_logic;
        in673 : in std_logic;
        in674 : in std_logic;
        in675 : in std_logic;
        in676 : in std_logic;
        in677 : in std_logic;
        in678 : in std_logic;
        in679 : in std_logic;
        in680 : in std_logic;
        in681 : in std_logic;
        in682 : in std_logic;
        in683 : in std_logic;
        in684 : in std_logic;
        in685 : in std_logic;
        in686 : in std_logic;
        in687 : in std_logic;
        in688 : in std_logic;
        in689 : in std_logic;
        in690 : in std_logic;
        in691 : in std_logic;
        in692 : in std_logic;
        in693 : in std_logic;
        in694 : in std_logic;
        in695 : in std_logic;
        in696 : in std_logic;
        in697 : in std_logic;
        in698 : in std_logic;
        in699 : in std_logic;
        in700 : in std_logic;
        in701 : in std_logic;
        in702 : in std_logic;
        in703 : in std_logic;
        in704 : in std_logic;
        in705 : in std_logic;
        in706 : in std_logic;
        in707 : in std_logic;
        in708 : in std_logic;
        in709 : in std_logic;
        in710 : in std_logic;
        in711 : in std_logic;
        in712 : in std_logic;
        in713 : in std_logic;
        in714 : in std_logic;
        in715 : in std_logic;
        in716 : in std_logic;
        in717 : in std_logic;
        in718 : in std_logic;
        in719 : in std_logic;
        in720 : in std_logic;
        in721 : in std_logic;
        in722 : in std_logic;
        in723 : in std_logic;
        in724 : in std_logic;
        in725 : in std_logic;
        in726 : in std_logic;
        in727 : in std_logic;
        in728 : in std_logic;
        in729 : in std_logic;
        in730 : in std_logic;
        in731 : in std_logic;
        in732 : in std_logic;
        in733 : in std_logic;
        in734 : in std_logic;
        in735 : in std_logic;
        in736 : in std_logic;
        in737 : in std_logic;
        in738 : in std_logic;
        in739 : in std_logic;
        in740 : in std_logic;
        in741 : in std_logic;
        in742 : in std_logic;
        in743 : in std_logic;
        in744 : in std_logic;
        in745 : in std_logic;
        in746 : in std_logic;
        in747 : in std_logic;
        in748 : in std_logic;
        in749 : in std_logic;
        in750 : in std_logic;
        in751 : in std_logic;
        in752 : in std_logic;
        in753 : in std_logic;
        in754 : in std_logic;
        in755 : in std_logic;
        in756 : in std_logic;
        in757 : in std_logic;
        in758 : in std_logic;
        in759 : in std_logic;
        in760 : in std_logic;
        in761 : in std_logic;
        in762 : in std_logic;
        in763 : in std_logic;
        in764 : in std_logic;
        in765 : in std_logic;
        in766 : in std_logic;
        in767 : in std_logic;
        in768 : in std_logic;
        in769 : in std_logic;
        in770 : in std_logic;
        in771 : in std_logic;
        in772 : in std_logic;
        in773 : in std_logic;
        in774 : in std_logic;
        in775 : in std_logic;
        in776 : in std_logic;
        in777 : in std_logic;
        in778 : in std_logic;
        in779 : in std_logic;
        in780 : in std_logic;
        in781 : in std_logic;
        in782 : in std_logic;
        in783 : in std_logic;
        in784 : in std_logic;
        in785 : in std_logic;
        in786 : in std_logic;
        in787 : in std_logic;
        in788 : in std_logic;
        in789 : in std_logic;
        in790 : in std_logic;
        in791 : in std_logic;
        in792 : in std_logic;
        in793 : in std_logic;
        in794 : in std_logic;
        in795 : in std_logic;
        in796 : in std_logic;
        in797 : in std_logic;
        in798 : in std_logic;
        in799 : in std_logic;
        in800 : in std_logic;
        in801 : in std_logic;
        in802 : in std_logic;
        in803 : in std_logic;
        in804 : in std_logic;
        in805 : in std_logic;
        in806 : in std_logic;
        in807 : in std_logic;
        in808 : in std_logic;
        in809 : in std_logic;
        in810 : in std_logic;
        in811 : in std_logic;
        in812 : in std_logic;
        in813 : in std_logic;
        in814 : in std_logic;
        in815 : in std_logic;
        in816 : in std_logic;
        in817 : in std_logic;
        in818 : in std_logic;
        in819 : in std_logic;
        in820 : in std_logic;
        in821 : in std_logic;
        in822 : in std_logic;
        in823 : in std_logic;
        in824 : in std_logic;
        in825 : in std_logic;
        in826 : in std_logic;
        in827 : in std_logic;
        in828 : in std_logic;
        in829 : in std_logic;
        in830 : in std_logic;
        in831 : in std_logic;
        in832 : in std_logic;
        in833 : in std_logic;
        in834 : in std_logic;
        in835 : in std_logic;
        in836 : in std_logic;
        in837 : in std_logic;
        in838 : in std_logic;
        in839 : in std_logic;
        in840 : in std_logic;
        in841 : in std_logic;
        in842 : in std_logic;
        in843 : in std_logic;
        in844 : in std_logic;
        in845 : in std_logic;
        in846 : in std_logic;
        in847 : in std_logic;
        in848 : in std_logic;
        in849 : in std_logic;
        in850 : in std_logic;
        in851 : in std_logic;
        in852 : in std_logic;
        in853 : in std_logic;
        in854 : in std_logic;
        in855 : in std_logic;
        in856 : in std_logic;
        in857 : in std_logic;
        in858 : in std_logic;
        in859 : in std_logic;
        in860 : in std_logic;
        in861 : in std_logic;
        in862 : in std_logic;
        in863 : in std_logic;
        in864 : in std_logic;
        in865 : in std_logic;
        in866 : in std_logic;
        in867 : in std_logic;
        in868 : in std_logic;
        in869 : in std_logic;
        in870 : in std_logic;
        in871 : in std_logic;
        in872 : in std_logic;
        in873 : in std_logic;
        in874 : in std_logic;
        in875 : in std_logic;
        in876 : in std_logic;
        in877 : in std_logic;
        in878 : in std_logic;
        in879 : in std_logic;
        in880 : in std_logic;
        in881 : in std_logic;
        in882 : in std_logic;
        in883 : in std_logic;
        in884 : in std_logic;
        in885 : in std_logic;
        in886 : in std_logic;
        in887 : in std_logic;
        in888 : in std_logic;
        in889 : in std_logic;
        in890 : in std_logic;
        in891 : in std_logic;
        in892 : in std_logic;
        in893 : in std_logic;
        in894 : in std_logic;
        in895 : in std_logic;
        in896 : in std_logic;
        in897 : in std_logic;
        in898 : in std_logic;
        in899 : in std_logic;
        in900 : in std_logic;
        in901 : in std_logic;
        in902 : in std_logic;
        in903 : in std_logic;
        in904 : in std_logic;
        in905 : in std_logic;
        in906 : in std_logic;
        in907 : in std_logic;
        in908 : in std_logic;
        in909 : in std_logic;
        in910 : in std_logic;
        in911 : in std_logic;
        in912 : in std_logic;
        in913 : in std_logic;
        in914 : in std_logic;
        in915 : in std_logic;
        in916 : in std_logic;
        in917 : in std_logic;
        in918 : in std_logic;
        in919 : in std_logic;
        in920 : in std_logic;
        in921 : in std_logic;
        in922 : in std_logic;
        in923 : in std_logic;
        in924 : in std_logic;
        in925 : in std_logic;
        in926 : in std_logic;
        in927 : in std_logic;
        in928 : in std_logic;
        in929 : in std_logic;
        in930 : in std_logic;
        in931 : in std_logic;
        in932 : in std_logic;
        in933 : in std_logic;
        in934 : in std_logic;
        in935 : in std_logic;
        in936 : in std_logic;
        in937 : in std_logic;
        in938 : in std_logic;
        in939 : in std_logic;
        in940 : in std_logic;
        in941 : in std_logic;
        in942 : in std_logic;
        in943 : in std_logic;
        in944 : in std_logic;
        in945 : in std_logic;
        in946 : in std_logic;
        in947 : in std_logic;
        in948 : in std_logic;
        in949 : in std_logic;
        in950 : in std_logic;
        in951 : in std_logic;
        in952 : in std_logic;
        in953 : in std_logic;
        in954 : in std_logic;
        in955 : in std_logic;
        in956 : in std_logic;
        in957 : in std_logic;
        in958 : in std_logic;
        in959 : in std_logic;
        in960 : in std_logic;
        in961 : in std_logic;
        in962 : in std_logic;
        in963 : in std_logic;
        in964 : in std_logic;
        in965 : in std_logic;
        in966 : in std_logic;
        in967 : in std_logic;
        in968 : in std_logic;
        in969 : in std_logic;
        in970 : in std_logic;
        in971 : in std_logic;
        in972 : in std_logic;
        in973 : in std_logic;
        in974 : in std_logic;
        in975 : in std_logic;
        in976 : in std_logic;
        in977 : in std_logic;
        in978 : in std_logic;
        in979 : in std_logic;
        in980 : in std_logic;
        in981 : in std_logic;
        in982 : in std_logic;
        in983 : in std_logic;
        in984 : in std_logic;
        in985 : in std_logic;
        in986 : in std_logic;
        in987 : in std_logic;
        in988 : in std_logic;
        in989 : in std_logic;
        in990 : in std_logic;
        in991 : in std_logic;
        in992 : in std_logic;
        in993 : in std_logic;
        in994 : in std_logic;
        in995 : in std_logic;
        in996 : in std_logic;
        in997 : in std_logic;
        in998 : in std_logic;
        in999 : in std_logic;
        in1000 : in std_logic;
        in1001 : in std_logic;
        in1002 : in std_logic;
        in1003 : in std_logic;
        in1004 : in std_logic;
        in1005 : in std_logic;
        in1006 : in std_logic;
        in1007 : in std_logic;
        in1008 : in std_logic;
        in1009 : in std_logic;
        in1010 : in std_logic;
        in1011 : in std_logic;
        in1012 : in std_logic;
        in1013 : in std_logic;
        in1014 : in std_logic;
        in1015 : in std_logic;
        in1016 : in std_logic;
        in1017 : in std_logic;
        in1018 : in std_logic;
        in1019 : in std_logic;
        in1020 : in std_logic;
        in1021 : in std_logic;
        in1022 : in std_logic;
        in1023 : in std_logic;
        mux_out : out std_logic
    );
end entity mux_1024to1;

architecture behavior of mux_1024to1 is


begin

    selection : process(mux_sel, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, in100, in101, in102, in103, in104, in105, in106, in107, in108, in109, in110, in111, in112, in113, in114, in115, in116, in117, in118, in119, in120, in121, in122, in123, in124, in125, in126, in127, in128, in129, in130, in131, in132, in133, in134, in135, in136, in137, in138, in139, in140, in141, in142, in143, in144, in145, in146, in147, in148, in149, in150, in151, in152, in153, in154, in155, in156, in157, in158, in159, in160, in161, in162, in163, in164, in165, in166, in167, in168, in169, in170, in171, in172, in173, in174, in175, in176, in177, in178, in179, in180, in181, in182, in183, in184, in185, in186, in187, in188, in189, in190, in191, in192, in193, in194, in195, in196, in197, in198, in199, in200, in201, in202, in203, in204, in205, in206, in207, in208, in209, in210, in211, in212, in213, in214, in215, in216, in217, in218, in219, in220, in221, in222, in223, in224, in225, in226, in227, in228, in229, in230, in231, in232, in233, in234, in235, in236, in237, in238, in239, in240, in241, in242, in243, in244, in245, in246, in247, in248, in249, in250, in251, in252, in253, in254, in255, in256, in257, in258, in259, in260, in261, in262, in263, in264, in265, in266, in267, in268, in269, in270, in271, in272, in273, in274, in275, in276, in277, in278, in279, in280, in281, in282, in283, in284, in285, in286, in287, in288, in289, in290, in291, in292, in293, in294, in295, in296, in297, in298, in299, in300, in301, in302, in303, in304, in305, in306, in307, in308, in309, in310, in311, in312, in313, in314, in315, in316, in317, in318, in319, in320, in321, in322, in323, in324, in325, in326, in327, in328, in329, in330, in331, in332, in333, in334, in335, in336, in337, in338, in339, in340, in341, in342, in343, in344, in345, in346, in347, in348, in349, in350, in351, in352, in353, in354, in355, in356, in357, in358, in359, in360, in361, in362, in363, in364, in365, in366, in367, in368, in369, in370, in371, in372, in373, in374, in375, in376, in377, in378, in379, in380, in381, in382, in383, in384, in385, in386, in387, in388, in389, in390, in391, in392, in393, in394, in395, in396, in397, in398, in399, in400, in401, in402, in403, in404, in405, in406, in407, in408, in409, in410, in411, in412, in413, in414, in415, in416, in417, in418, in419, in420, in421, in422, in423, in424, in425, in426, in427, in428, in429, in430, in431, in432, in433, in434, in435, in436, in437, in438, in439, in440, in441, in442, in443, in444, in445, in446, in447, in448, in449, in450, in451, in452, in453, in454, in455, in456, in457, in458, in459, in460, in461, in462, in463, in464, in465, in466, in467, in468, in469, in470, in471, in472, in473, in474, in475, in476, in477, in478, in479, in480, in481, in482, in483, in484, in485, in486, in487, in488, in489, in490, in491, in492, in493, in494, in495, in496, in497, in498, in499, in500, in501, in502, in503, in504, in505, in506, in507, in508, in509, in510, in511, in512, in513, in514, in515, in516, in517, in518, in519, in520, in521, in522, in523, in524, in525, in526, in527, in528, in529, in530, in531, in532, in533, in534, in535, in536, in537, in538, in539, in540, in541, in542, in543, in544, in545, in546, in547, in548, in549, in550, in551, in552, in553, in554, in555, in556, in557, in558, in559, in560, in561, in562, in563, in564, in565, in566, in567, in568, in569, in570, in571, in572, in573, in574, in575, in576, in577, in578, in579, in580, in581, in582, in583, in584, in585, in586, in587, in588, in589, in590, in591, in592, in593, in594, in595, in596, in597, in598, in599, in600, in601, in602, in603, in604, in605, in606, in607, in608, in609, in610, in611, in612, in613, in614, in615, in616, in617, in618, in619, in620, in621, in622, in623, in624, in625, in626, in627, in628, in629, in630, in631, in632, in633, in634, in635, in636, in637, in638, in639, in640, in641, in642, in643, in644, in645, in646, in647, in648, in649, in650, in651, in652, in653, in654, in655, in656, in657, in658, in659, in660, in661, in662, in663, in664, in665, in666, in667, in668, in669, in670, in671, in672, in673, in674, in675, in676, in677, in678, in679, in680, in681, in682, in683, in684, in685, in686, in687, in688, in689, in690, in691, in692, in693, in694, in695, in696, in697, in698, in699, in700, in701, in702, in703, in704, in705, in706, in707, in708, in709, in710, in711, in712, in713, in714, in715, in716, in717, in718, in719, in720, in721, in722, in723, in724, in725, in726, in727, in728, in729, in730, in731, in732, in733, in734, in735, in736, in737, in738, in739, in740, in741, in742, in743, in744, in745, in746, in747, in748, in749, in750, in751, in752, in753, in754, in755, in756, in757, in758, in759, in760, in761, in762, in763, in764, in765, in766, in767, in768, in769, in770, in771, in772, in773, in774, in775, in776, in777, in778, in779, in780, in781, in782, in783, in784, in785, in786, in787, in788, in789, in790, in791, in792, in793, in794, in795, in796, in797, in798, in799, in800, in801, in802, in803, in804, in805, in806, in807, in808, in809, in810, in811, in812, in813, in814, in815, in816, in817, in818, in819, in820, in821, in822, in823, in824, in825, in826, in827, in828, in829, in830, in831, in832, in833, in834, in835, in836, in837, in838, in839, in840, in841, in842, in843, in844, in845, in846, in847, in848, in849, in850, in851, in852, in853, in854, in855, in856, in857, in858, in859, in860, in861, in862, in863, in864, in865, in866, in867, in868, in869, in870, in871, in872, in873, in874, in875, in876, in877, in878, in879, in880, in881, in882, in883, in884, in885, in886, in887, in888, in889, in890, in891, in892, in893, in894, in895, in896, in897, in898, in899, in900, in901, in902, in903, in904, in905, in906, in907, in908, in909, in910, in911, in912, in913, in914, in915, in916, in917, in918, in919, in920, in921, in922, in923, in924, in925, in926, in927, in928, in929, in930, in931, in932, in933, in934, in935, in936, in937, in938, in939, in940, in941, in942, in943, in944, in945, in946, in947, in948, in949, in950, in951, in952, in953, in954, in955, in956, in957, in958, in959, in960, in961, in962, in963, in964, in965, in966, in967, in968, in969, in970, in971, in972, in973, in974, in975, in976, in977, in978, in979, in980, in981, in982, in983, in984, in985, in986, in987, in988, in989, in990, in991, in992, in993, in994, in995, in996, in997, in998, in999, in1000, in1001, in1002, in1003, in1004, in1005, in1006, in1007, in1008, in1009, in1010, in1011, in1012, in1013, in1014, in1015, in1016, in1017, in1018, in1019, in1020, in1021, in1022, in1023 )
    begin

        case mux_sel is

            when "0000000000" =>
                mux_out <= in0;


            when "0000000001" =>
                mux_out <= in1;


            when "0000000010" =>
                mux_out <= in2;


            when "0000000011" =>
                mux_out <= in3;


            when "0000000100" =>
                mux_out <= in4;


            when "0000000101" =>
                mux_out <= in5;


            when "0000000110" =>
                mux_out <= in6;


            when "0000000111" =>
                mux_out <= in7;


            when "0000001000" =>
                mux_out <= in8;


            when "0000001001" =>
                mux_out <= in9;


            when "0000001010" =>
                mux_out <= in10;


            when "0000001011" =>
                mux_out <= in11;


            when "0000001100" =>
                mux_out <= in12;


            when "0000001101" =>
                mux_out <= in13;


            when "0000001110" =>
                mux_out <= in14;


            when "0000001111" =>
                mux_out <= in15;


            when "0000010000" =>
                mux_out <= in16;


            when "0000010001" =>
                mux_out <= in17;


            when "0000010010" =>
                mux_out <= in18;


            when "0000010011" =>
                mux_out <= in19;


            when "0000010100" =>
                mux_out <= in20;


            when "0000010101" =>
                mux_out <= in21;


            when "0000010110" =>
                mux_out <= in22;


            when "0000010111" =>
                mux_out <= in23;


            when "0000011000" =>
                mux_out <= in24;


            when "0000011001" =>
                mux_out <= in25;


            when "0000011010" =>
                mux_out <= in26;


            when "0000011011" =>
                mux_out <= in27;


            when "0000011100" =>
                mux_out <= in28;


            when "0000011101" =>
                mux_out <= in29;


            when "0000011110" =>
                mux_out <= in30;


            when "0000011111" =>
                mux_out <= in31;


            when "0000100000" =>
                mux_out <= in32;


            when "0000100001" =>
                mux_out <= in33;


            when "0000100010" =>
                mux_out <= in34;


            when "0000100011" =>
                mux_out <= in35;


            when "0000100100" =>
                mux_out <= in36;


            when "0000100101" =>
                mux_out <= in37;


            when "0000100110" =>
                mux_out <= in38;


            when "0000100111" =>
                mux_out <= in39;


            when "0000101000" =>
                mux_out <= in40;


            when "0000101001" =>
                mux_out <= in41;


            when "0000101010" =>
                mux_out <= in42;


            when "0000101011" =>
                mux_out <= in43;


            when "0000101100" =>
                mux_out <= in44;


            when "0000101101" =>
                mux_out <= in45;


            when "0000101110" =>
                mux_out <= in46;


            when "0000101111" =>
                mux_out <= in47;


            when "0000110000" =>
                mux_out <= in48;


            when "0000110001" =>
                mux_out <= in49;


            when "0000110010" =>
                mux_out <= in50;


            when "0000110011" =>
                mux_out <= in51;


            when "0000110100" =>
                mux_out <= in52;


            when "0000110101" =>
                mux_out <= in53;


            when "0000110110" =>
                mux_out <= in54;


            when "0000110111" =>
                mux_out <= in55;


            when "0000111000" =>
                mux_out <= in56;


            when "0000111001" =>
                mux_out <= in57;


            when "0000111010" =>
                mux_out <= in58;


            when "0000111011" =>
                mux_out <= in59;


            when "0000111100" =>
                mux_out <= in60;


            when "0000111101" =>
                mux_out <= in61;


            when "0000111110" =>
                mux_out <= in62;


            when "0000111111" =>
                mux_out <= in63;


            when "0001000000" =>
                mux_out <= in64;


            when "0001000001" =>
                mux_out <= in65;


            when "0001000010" =>
                mux_out <= in66;


            when "0001000011" =>
                mux_out <= in67;


            when "0001000100" =>
                mux_out <= in68;


            when "0001000101" =>
                mux_out <= in69;


            when "0001000110" =>
                mux_out <= in70;


            when "0001000111" =>
                mux_out <= in71;


            when "0001001000" =>
                mux_out <= in72;


            when "0001001001" =>
                mux_out <= in73;


            when "0001001010" =>
                mux_out <= in74;


            when "0001001011" =>
                mux_out <= in75;


            when "0001001100" =>
                mux_out <= in76;


            when "0001001101" =>
                mux_out <= in77;


            when "0001001110" =>
                mux_out <= in78;


            when "0001001111" =>
                mux_out <= in79;


            when "0001010000" =>
                mux_out <= in80;


            when "0001010001" =>
                mux_out <= in81;


            when "0001010010" =>
                mux_out <= in82;


            when "0001010011" =>
                mux_out <= in83;


            when "0001010100" =>
                mux_out <= in84;


            when "0001010101" =>
                mux_out <= in85;


            when "0001010110" =>
                mux_out <= in86;


            when "0001010111" =>
                mux_out <= in87;


            when "0001011000" =>
                mux_out <= in88;


            when "0001011001" =>
                mux_out <= in89;


            when "0001011010" =>
                mux_out <= in90;


            when "0001011011" =>
                mux_out <= in91;


            when "0001011100" =>
                mux_out <= in92;


            when "0001011101" =>
                mux_out <= in93;


            when "0001011110" =>
                mux_out <= in94;


            when "0001011111" =>
                mux_out <= in95;


            when "0001100000" =>
                mux_out <= in96;


            when "0001100001" =>
                mux_out <= in97;


            when "0001100010" =>
                mux_out <= in98;


            when "0001100011" =>
                mux_out <= in99;


            when "0001100100" =>
                mux_out <= in100;


            when "0001100101" =>
                mux_out <= in101;


            when "0001100110" =>
                mux_out <= in102;


            when "0001100111" =>
                mux_out <= in103;


            when "0001101000" =>
                mux_out <= in104;


            when "0001101001" =>
                mux_out <= in105;


            when "0001101010" =>
                mux_out <= in106;


            when "0001101011" =>
                mux_out <= in107;


            when "0001101100" =>
                mux_out <= in108;


            when "0001101101" =>
                mux_out <= in109;


            when "0001101110" =>
                mux_out <= in110;


            when "0001101111" =>
                mux_out <= in111;


            when "0001110000" =>
                mux_out <= in112;


            when "0001110001" =>
                mux_out <= in113;


            when "0001110010" =>
                mux_out <= in114;


            when "0001110011" =>
                mux_out <= in115;


            when "0001110100" =>
                mux_out <= in116;


            when "0001110101" =>
                mux_out <= in117;


            when "0001110110" =>
                mux_out <= in118;


            when "0001110111" =>
                mux_out <= in119;


            when "0001111000" =>
                mux_out <= in120;


            when "0001111001" =>
                mux_out <= in121;


            when "0001111010" =>
                mux_out <= in122;


            when "0001111011" =>
                mux_out <= in123;


            when "0001111100" =>
                mux_out <= in124;


            when "0001111101" =>
                mux_out <= in125;


            when "0001111110" =>
                mux_out <= in126;


            when "0001111111" =>
                mux_out <= in127;


            when "0010000000" =>
                mux_out <= in128;


            when "0010000001" =>
                mux_out <= in129;


            when "0010000010" =>
                mux_out <= in130;


            when "0010000011" =>
                mux_out <= in131;


            when "0010000100" =>
                mux_out <= in132;


            when "0010000101" =>
                mux_out <= in133;


            when "0010000110" =>
                mux_out <= in134;


            when "0010000111" =>
                mux_out <= in135;


            when "0010001000" =>
                mux_out <= in136;


            when "0010001001" =>
                mux_out <= in137;


            when "0010001010" =>
                mux_out <= in138;


            when "0010001011" =>
                mux_out <= in139;


            when "0010001100" =>
                mux_out <= in140;


            when "0010001101" =>
                mux_out <= in141;


            when "0010001110" =>
                mux_out <= in142;


            when "0010001111" =>
                mux_out <= in143;


            when "0010010000" =>
                mux_out <= in144;


            when "0010010001" =>
                mux_out <= in145;


            when "0010010010" =>
                mux_out <= in146;


            when "0010010011" =>
                mux_out <= in147;


            when "0010010100" =>
                mux_out <= in148;


            when "0010010101" =>
                mux_out <= in149;


            when "0010010110" =>
                mux_out <= in150;


            when "0010010111" =>
                mux_out <= in151;


            when "0010011000" =>
                mux_out <= in152;


            when "0010011001" =>
                mux_out <= in153;


            when "0010011010" =>
                mux_out <= in154;


            when "0010011011" =>
                mux_out <= in155;


            when "0010011100" =>
                mux_out <= in156;


            when "0010011101" =>
                mux_out <= in157;


            when "0010011110" =>
                mux_out <= in158;


            when "0010011111" =>
                mux_out <= in159;


            when "0010100000" =>
                mux_out <= in160;


            when "0010100001" =>
                mux_out <= in161;


            when "0010100010" =>
                mux_out <= in162;


            when "0010100011" =>
                mux_out <= in163;


            when "0010100100" =>
                mux_out <= in164;


            when "0010100101" =>
                mux_out <= in165;


            when "0010100110" =>
                mux_out <= in166;


            when "0010100111" =>
                mux_out <= in167;


            when "0010101000" =>
                mux_out <= in168;


            when "0010101001" =>
                mux_out <= in169;


            when "0010101010" =>
                mux_out <= in170;


            when "0010101011" =>
                mux_out <= in171;


            when "0010101100" =>
                mux_out <= in172;


            when "0010101101" =>
                mux_out <= in173;


            when "0010101110" =>
                mux_out <= in174;


            when "0010101111" =>
                mux_out <= in175;


            when "0010110000" =>
                mux_out <= in176;


            when "0010110001" =>
                mux_out <= in177;


            when "0010110010" =>
                mux_out <= in178;


            when "0010110011" =>
                mux_out <= in179;


            when "0010110100" =>
                mux_out <= in180;


            when "0010110101" =>
                mux_out <= in181;


            when "0010110110" =>
                mux_out <= in182;


            when "0010110111" =>
                mux_out <= in183;


            when "0010111000" =>
                mux_out <= in184;


            when "0010111001" =>
                mux_out <= in185;


            when "0010111010" =>
                mux_out <= in186;


            when "0010111011" =>
                mux_out <= in187;


            when "0010111100" =>
                mux_out <= in188;


            when "0010111101" =>
                mux_out <= in189;


            when "0010111110" =>
                mux_out <= in190;


            when "0010111111" =>
                mux_out <= in191;


            when "0011000000" =>
                mux_out <= in192;


            when "0011000001" =>
                mux_out <= in193;


            when "0011000010" =>
                mux_out <= in194;


            when "0011000011" =>
                mux_out <= in195;


            when "0011000100" =>
                mux_out <= in196;


            when "0011000101" =>
                mux_out <= in197;


            when "0011000110" =>
                mux_out <= in198;


            when "0011000111" =>
                mux_out <= in199;


            when "0011001000" =>
                mux_out <= in200;


            when "0011001001" =>
                mux_out <= in201;


            when "0011001010" =>
                mux_out <= in202;


            when "0011001011" =>
                mux_out <= in203;


            when "0011001100" =>
                mux_out <= in204;


            when "0011001101" =>
                mux_out <= in205;


            when "0011001110" =>
                mux_out <= in206;


            when "0011001111" =>
                mux_out <= in207;


            when "0011010000" =>
                mux_out <= in208;


            when "0011010001" =>
                mux_out <= in209;


            when "0011010010" =>
                mux_out <= in210;


            when "0011010011" =>
                mux_out <= in211;


            when "0011010100" =>
                mux_out <= in212;


            when "0011010101" =>
                mux_out <= in213;


            when "0011010110" =>
                mux_out <= in214;


            when "0011010111" =>
                mux_out <= in215;


            when "0011011000" =>
                mux_out <= in216;


            when "0011011001" =>
                mux_out <= in217;


            when "0011011010" =>
                mux_out <= in218;


            when "0011011011" =>
                mux_out <= in219;


            when "0011011100" =>
                mux_out <= in220;


            when "0011011101" =>
                mux_out <= in221;


            when "0011011110" =>
                mux_out <= in222;


            when "0011011111" =>
                mux_out <= in223;


            when "0011100000" =>
                mux_out <= in224;


            when "0011100001" =>
                mux_out <= in225;


            when "0011100010" =>
                mux_out <= in226;


            when "0011100011" =>
                mux_out <= in227;


            when "0011100100" =>
                mux_out <= in228;


            when "0011100101" =>
                mux_out <= in229;


            when "0011100110" =>
                mux_out <= in230;


            when "0011100111" =>
                mux_out <= in231;


            when "0011101000" =>
                mux_out <= in232;


            when "0011101001" =>
                mux_out <= in233;


            when "0011101010" =>
                mux_out <= in234;


            when "0011101011" =>
                mux_out <= in235;


            when "0011101100" =>
                mux_out <= in236;


            when "0011101101" =>
                mux_out <= in237;


            when "0011101110" =>
                mux_out <= in238;


            when "0011101111" =>
                mux_out <= in239;


            when "0011110000" =>
                mux_out <= in240;


            when "0011110001" =>
                mux_out <= in241;


            when "0011110010" =>
                mux_out <= in242;


            when "0011110011" =>
                mux_out <= in243;


            when "0011110100" =>
                mux_out <= in244;


            when "0011110101" =>
                mux_out <= in245;


            when "0011110110" =>
                mux_out <= in246;


            when "0011110111" =>
                mux_out <= in247;


            when "0011111000" =>
                mux_out <= in248;


            when "0011111001" =>
                mux_out <= in249;


            when "0011111010" =>
                mux_out <= in250;


            when "0011111011" =>
                mux_out <= in251;


            when "0011111100" =>
                mux_out <= in252;


            when "0011111101" =>
                mux_out <= in253;


            when "0011111110" =>
                mux_out <= in254;


            when "0011111111" =>
                mux_out <= in255;


            when "0100000000" =>
                mux_out <= in256;


            when "0100000001" =>
                mux_out <= in257;


            when "0100000010" =>
                mux_out <= in258;


            when "0100000011" =>
                mux_out <= in259;


            when "0100000100" =>
                mux_out <= in260;


            when "0100000101" =>
                mux_out <= in261;


            when "0100000110" =>
                mux_out <= in262;


            when "0100000111" =>
                mux_out <= in263;


            when "0100001000" =>
                mux_out <= in264;


            when "0100001001" =>
                mux_out <= in265;


            when "0100001010" =>
                mux_out <= in266;


            when "0100001011" =>
                mux_out <= in267;


            when "0100001100" =>
                mux_out <= in268;


            when "0100001101" =>
                mux_out <= in269;


            when "0100001110" =>
                mux_out <= in270;


            when "0100001111" =>
                mux_out <= in271;


            when "0100010000" =>
                mux_out <= in272;


            when "0100010001" =>
                mux_out <= in273;


            when "0100010010" =>
                mux_out <= in274;


            when "0100010011" =>
                mux_out <= in275;


            when "0100010100" =>
                mux_out <= in276;


            when "0100010101" =>
                mux_out <= in277;


            when "0100010110" =>
                mux_out <= in278;


            when "0100010111" =>
                mux_out <= in279;


            when "0100011000" =>
                mux_out <= in280;


            when "0100011001" =>
                mux_out <= in281;


            when "0100011010" =>
                mux_out <= in282;


            when "0100011011" =>
                mux_out <= in283;


            when "0100011100" =>
                mux_out <= in284;


            when "0100011101" =>
                mux_out <= in285;


            when "0100011110" =>
                mux_out <= in286;


            when "0100011111" =>
                mux_out <= in287;


            when "0100100000" =>
                mux_out <= in288;


            when "0100100001" =>
                mux_out <= in289;


            when "0100100010" =>
                mux_out <= in290;


            when "0100100011" =>
                mux_out <= in291;


            when "0100100100" =>
                mux_out <= in292;


            when "0100100101" =>
                mux_out <= in293;


            when "0100100110" =>
                mux_out <= in294;


            when "0100100111" =>
                mux_out <= in295;


            when "0100101000" =>
                mux_out <= in296;


            when "0100101001" =>
                mux_out <= in297;


            when "0100101010" =>
                mux_out <= in298;


            when "0100101011" =>
                mux_out <= in299;


            when "0100101100" =>
                mux_out <= in300;


            when "0100101101" =>
                mux_out <= in301;


            when "0100101110" =>
                mux_out <= in302;


            when "0100101111" =>
                mux_out <= in303;


            when "0100110000" =>
                mux_out <= in304;


            when "0100110001" =>
                mux_out <= in305;


            when "0100110010" =>
                mux_out <= in306;


            when "0100110011" =>
                mux_out <= in307;


            when "0100110100" =>
                mux_out <= in308;


            when "0100110101" =>
                mux_out <= in309;


            when "0100110110" =>
                mux_out <= in310;


            when "0100110111" =>
                mux_out <= in311;


            when "0100111000" =>
                mux_out <= in312;


            when "0100111001" =>
                mux_out <= in313;


            when "0100111010" =>
                mux_out <= in314;


            when "0100111011" =>
                mux_out <= in315;


            when "0100111100" =>
                mux_out <= in316;


            when "0100111101" =>
                mux_out <= in317;


            when "0100111110" =>
                mux_out <= in318;


            when "0100111111" =>
                mux_out <= in319;


            when "0101000000" =>
                mux_out <= in320;


            when "0101000001" =>
                mux_out <= in321;


            when "0101000010" =>
                mux_out <= in322;


            when "0101000011" =>
                mux_out <= in323;


            when "0101000100" =>
                mux_out <= in324;


            when "0101000101" =>
                mux_out <= in325;


            when "0101000110" =>
                mux_out <= in326;


            when "0101000111" =>
                mux_out <= in327;


            when "0101001000" =>
                mux_out <= in328;


            when "0101001001" =>
                mux_out <= in329;


            when "0101001010" =>
                mux_out <= in330;


            when "0101001011" =>
                mux_out <= in331;


            when "0101001100" =>
                mux_out <= in332;


            when "0101001101" =>
                mux_out <= in333;


            when "0101001110" =>
                mux_out <= in334;


            when "0101001111" =>
                mux_out <= in335;


            when "0101010000" =>
                mux_out <= in336;


            when "0101010001" =>
                mux_out <= in337;


            when "0101010010" =>
                mux_out <= in338;


            when "0101010011" =>
                mux_out <= in339;


            when "0101010100" =>
                mux_out <= in340;


            when "0101010101" =>
                mux_out <= in341;


            when "0101010110" =>
                mux_out <= in342;


            when "0101010111" =>
                mux_out <= in343;


            when "0101011000" =>
                mux_out <= in344;


            when "0101011001" =>
                mux_out <= in345;


            when "0101011010" =>
                mux_out <= in346;


            when "0101011011" =>
                mux_out <= in347;


            when "0101011100" =>
                mux_out <= in348;


            when "0101011101" =>
                mux_out <= in349;


            when "0101011110" =>
                mux_out <= in350;


            when "0101011111" =>
                mux_out <= in351;


            when "0101100000" =>
                mux_out <= in352;


            when "0101100001" =>
                mux_out <= in353;


            when "0101100010" =>
                mux_out <= in354;


            when "0101100011" =>
                mux_out <= in355;


            when "0101100100" =>
                mux_out <= in356;


            when "0101100101" =>
                mux_out <= in357;


            when "0101100110" =>
                mux_out <= in358;


            when "0101100111" =>
                mux_out <= in359;


            when "0101101000" =>
                mux_out <= in360;


            when "0101101001" =>
                mux_out <= in361;


            when "0101101010" =>
                mux_out <= in362;


            when "0101101011" =>
                mux_out <= in363;


            when "0101101100" =>
                mux_out <= in364;


            when "0101101101" =>
                mux_out <= in365;


            when "0101101110" =>
                mux_out <= in366;


            when "0101101111" =>
                mux_out <= in367;


            when "0101110000" =>
                mux_out <= in368;


            when "0101110001" =>
                mux_out <= in369;


            when "0101110010" =>
                mux_out <= in370;


            when "0101110011" =>
                mux_out <= in371;


            when "0101110100" =>
                mux_out <= in372;


            when "0101110101" =>
                mux_out <= in373;


            when "0101110110" =>
                mux_out <= in374;


            when "0101110111" =>
                mux_out <= in375;


            when "0101111000" =>
                mux_out <= in376;


            when "0101111001" =>
                mux_out <= in377;


            when "0101111010" =>
                mux_out <= in378;


            when "0101111011" =>
                mux_out <= in379;


            when "0101111100" =>
                mux_out <= in380;


            when "0101111101" =>
                mux_out <= in381;


            when "0101111110" =>
                mux_out <= in382;


            when "0101111111" =>
                mux_out <= in383;


            when "0110000000" =>
                mux_out <= in384;


            when "0110000001" =>
                mux_out <= in385;


            when "0110000010" =>
                mux_out <= in386;


            when "0110000011" =>
                mux_out <= in387;


            when "0110000100" =>
                mux_out <= in388;


            when "0110000101" =>
                mux_out <= in389;


            when "0110000110" =>
                mux_out <= in390;


            when "0110000111" =>
                mux_out <= in391;


            when "0110001000" =>
                mux_out <= in392;


            when "0110001001" =>
                mux_out <= in393;


            when "0110001010" =>
                mux_out <= in394;


            when "0110001011" =>
                mux_out <= in395;


            when "0110001100" =>
                mux_out <= in396;


            when "0110001101" =>
                mux_out <= in397;


            when "0110001110" =>
                mux_out <= in398;


            when "0110001111" =>
                mux_out <= in399;


            when "0110010000" =>
                mux_out <= in400;


            when "0110010001" =>
                mux_out <= in401;


            when "0110010010" =>
                mux_out <= in402;


            when "0110010011" =>
                mux_out <= in403;


            when "0110010100" =>
                mux_out <= in404;


            when "0110010101" =>
                mux_out <= in405;


            when "0110010110" =>
                mux_out <= in406;


            when "0110010111" =>
                mux_out <= in407;


            when "0110011000" =>
                mux_out <= in408;


            when "0110011001" =>
                mux_out <= in409;


            when "0110011010" =>
                mux_out <= in410;


            when "0110011011" =>
                mux_out <= in411;


            when "0110011100" =>
                mux_out <= in412;


            when "0110011101" =>
                mux_out <= in413;


            when "0110011110" =>
                mux_out <= in414;


            when "0110011111" =>
                mux_out <= in415;


            when "0110100000" =>
                mux_out <= in416;


            when "0110100001" =>
                mux_out <= in417;


            when "0110100010" =>
                mux_out <= in418;


            when "0110100011" =>
                mux_out <= in419;


            when "0110100100" =>
                mux_out <= in420;


            when "0110100101" =>
                mux_out <= in421;


            when "0110100110" =>
                mux_out <= in422;


            when "0110100111" =>
                mux_out <= in423;


            when "0110101000" =>
                mux_out <= in424;


            when "0110101001" =>
                mux_out <= in425;


            when "0110101010" =>
                mux_out <= in426;


            when "0110101011" =>
                mux_out <= in427;


            when "0110101100" =>
                mux_out <= in428;


            when "0110101101" =>
                mux_out <= in429;


            when "0110101110" =>
                mux_out <= in430;


            when "0110101111" =>
                mux_out <= in431;


            when "0110110000" =>
                mux_out <= in432;


            when "0110110001" =>
                mux_out <= in433;


            when "0110110010" =>
                mux_out <= in434;


            when "0110110011" =>
                mux_out <= in435;


            when "0110110100" =>
                mux_out <= in436;


            when "0110110101" =>
                mux_out <= in437;


            when "0110110110" =>
                mux_out <= in438;


            when "0110110111" =>
                mux_out <= in439;


            when "0110111000" =>
                mux_out <= in440;


            when "0110111001" =>
                mux_out <= in441;


            when "0110111010" =>
                mux_out <= in442;


            when "0110111011" =>
                mux_out <= in443;


            when "0110111100" =>
                mux_out <= in444;


            when "0110111101" =>
                mux_out <= in445;


            when "0110111110" =>
                mux_out <= in446;


            when "0110111111" =>
                mux_out <= in447;


            when "0111000000" =>
                mux_out <= in448;


            when "0111000001" =>
                mux_out <= in449;


            when "0111000010" =>
                mux_out <= in450;


            when "0111000011" =>
                mux_out <= in451;


            when "0111000100" =>
                mux_out <= in452;


            when "0111000101" =>
                mux_out <= in453;


            when "0111000110" =>
                mux_out <= in454;


            when "0111000111" =>
                mux_out <= in455;


            when "0111001000" =>
                mux_out <= in456;


            when "0111001001" =>
                mux_out <= in457;


            when "0111001010" =>
                mux_out <= in458;


            when "0111001011" =>
                mux_out <= in459;


            when "0111001100" =>
                mux_out <= in460;


            when "0111001101" =>
                mux_out <= in461;


            when "0111001110" =>
                mux_out <= in462;


            when "0111001111" =>
                mux_out <= in463;


            when "0111010000" =>
                mux_out <= in464;


            when "0111010001" =>
                mux_out <= in465;


            when "0111010010" =>
                mux_out <= in466;


            when "0111010011" =>
                mux_out <= in467;


            when "0111010100" =>
                mux_out <= in468;


            when "0111010101" =>
                mux_out <= in469;


            when "0111010110" =>
                mux_out <= in470;


            when "0111010111" =>
                mux_out <= in471;


            when "0111011000" =>
                mux_out <= in472;


            when "0111011001" =>
                mux_out <= in473;


            when "0111011010" =>
                mux_out <= in474;


            when "0111011011" =>
                mux_out <= in475;


            when "0111011100" =>
                mux_out <= in476;


            when "0111011101" =>
                mux_out <= in477;


            when "0111011110" =>
                mux_out <= in478;


            when "0111011111" =>
                mux_out <= in479;


            when "0111100000" =>
                mux_out <= in480;


            when "0111100001" =>
                mux_out <= in481;


            when "0111100010" =>
                mux_out <= in482;


            when "0111100011" =>
                mux_out <= in483;


            when "0111100100" =>
                mux_out <= in484;


            when "0111100101" =>
                mux_out <= in485;


            when "0111100110" =>
                mux_out <= in486;


            when "0111100111" =>
                mux_out <= in487;


            when "0111101000" =>
                mux_out <= in488;


            when "0111101001" =>
                mux_out <= in489;


            when "0111101010" =>
                mux_out <= in490;


            when "0111101011" =>
                mux_out <= in491;


            when "0111101100" =>
                mux_out <= in492;


            when "0111101101" =>
                mux_out <= in493;


            when "0111101110" =>
                mux_out <= in494;


            when "0111101111" =>
                mux_out <= in495;


            when "0111110000" =>
                mux_out <= in496;


            when "0111110001" =>
                mux_out <= in497;


            when "0111110010" =>
                mux_out <= in498;


            when "0111110011" =>
                mux_out <= in499;


            when "0111110100" =>
                mux_out <= in500;


            when "0111110101" =>
                mux_out <= in501;


            when "0111110110" =>
                mux_out <= in502;


            when "0111110111" =>
                mux_out <= in503;


            when "0111111000" =>
                mux_out <= in504;


            when "0111111001" =>
                mux_out <= in505;


            when "0111111010" =>
                mux_out <= in506;


            when "0111111011" =>
                mux_out <= in507;


            when "0111111100" =>
                mux_out <= in508;


            when "0111111101" =>
                mux_out <= in509;


            when "0111111110" =>
                mux_out <= in510;


            when "0111111111" =>
                mux_out <= in511;


            when "1000000000" =>
                mux_out <= in512;


            when "1000000001" =>
                mux_out <= in513;


            when "1000000010" =>
                mux_out <= in514;


            when "1000000011" =>
                mux_out <= in515;


            when "1000000100" =>
                mux_out <= in516;


            when "1000000101" =>
                mux_out <= in517;


            when "1000000110" =>
                mux_out <= in518;


            when "1000000111" =>
                mux_out <= in519;


            when "1000001000" =>
                mux_out <= in520;


            when "1000001001" =>
                mux_out <= in521;


            when "1000001010" =>
                mux_out <= in522;


            when "1000001011" =>
                mux_out <= in523;


            when "1000001100" =>
                mux_out <= in524;


            when "1000001101" =>
                mux_out <= in525;


            when "1000001110" =>
                mux_out <= in526;


            when "1000001111" =>
                mux_out <= in527;


            when "1000010000" =>
                mux_out <= in528;


            when "1000010001" =>
                mux_out <= in529;


            when "1000010010" =>
                mux_out <= in530;


            when "1000010011" =>
                mux_out <= in531;


            when "1000010100" =>
                mux_out <= in532;


            when "1000010101" =>
                mux_out <= in533;


            when "1000010110" =>
                mux_out <= in534;


            when "1000010111" =>
                mux_out <= in535;


            when "1000011000" =>
                mux_out <= in536;


            when "1000011001" =>
                mux_out <= in537;


            when "1000011010" =>
                mux_out <= in538;


            when "1000011011" =>
                mux_out <= in539;


            when "1000011100" =>
                mux_out <= in540;


            when "1000011101" =>
                mux_out <= in541;


            when "1000011110" =>
                mux_out <= in542;


            when "1000011111" =>
                mux_out <= in543;


            when "1000100000" =>
                mux_out <= in544;


            when "1000100001" =>
                mux_out <= in545;


            when "1000100010" =>
                mux_out <= in546;


            when "1000100011" =>
                mux_out <= in547;


            when "1000100100" =>
                mux_out <= in548;


            when "1000100101" =>
                mux_out <= in549;


            when "1000100110" =>
                mux_out <= in550;


            when "1000100111" =>
                mux_out <= in551;


            when "1000101000" =>
                mux_out <= in552;


            when "1000101001" =>
                mux_out <= in553;


            when "1000101010" =>
                mux_out <= in554;


            when "1000101011" =>
                mux_out <= in555;


            when "1000101100" =>
                mux_out <= in556;


            when "1000101101" =>
                mux_out <= in557;


            when "1000101110" =>
                mux_out <= in558;


            when "1000101111" =>
                mux_out <= in559;


            when "1000110000" =>
                mux_out <= in560;


            when "1000110001" =>
                mux_out <= in561;


            when "1000110010" =>
                mux_out <= in562;


            when "1000110011" =>
                mux_out <= in563;


            when "1000110100" =>
                mux_out <= in564;


            when "1000110101" =>
                mux_out <= in565;


            when "1000110110" =>
                mux_out <= in566;


            when "1000110111" =>
                mux_out <= in567;


            when "1000111000" =>
                mux_out <= in568;


            when "1000111001" =>
                mux_out <= in569;


            when "1000111010" =>
                mux_out <= in570;


            when "1000111011" =>
                mux_out <= in571;


            when "1000111100" =>
                mux_out <= in572;


            when "1000111101" =>
                mux_out <= in573;


            when "1000111110" =>
                mux_out <= in574;


            when "1000111111" =>
                mux_out <= in575;


            when "1001000000" =>
                mux_out <= in576;


            when "1001000001" =>
                mux_out <= in577;


            when "1001000010" =>
                mux_out <= in578;


            when "1001000011" =>
                mux_out <= in579;


            when "1001000100" =>
                mux_out <= in580;


            when "1001000101" =>
                mux_out <= in581;


            when "1001000110" =>
                mux_out <= in582;


            when "1001000111" =>
                mux_out <= in583;


            when "1001001000" =>
                mux_out <= in584;


            when "1001001001" =>
                mux_out <= in585;


            when "1001001010" =>
                mux_out <= in586;


            when "1001001011" =>
                mux_out <= in587;


            when "1001001100" =>
                mux_out <= in588;


            when "1001001101" =>
                mux_out <= in589;


            when "1001001110" =>
                mux_out <= in590;


            when "1001001111" =>
                mux_out <= in591;


            when "1001010000" =>
                mux_out <= in592;


            when "1001010001" =>
                mux_out <= in593;


            when "1001010010" =>
                mux_out <= in594;


            when "1001010011" =>
                mux_out <= in595;


            when "1001010100" =>
                mux_out <= in596;


            when "1001010101" =>
                mux_out <= in597;


            when "1001010110" =>
                mux_out <= in598;


            when "1001010111" =>
                mux_out <= in599;


            when "1001011000" =>
                mux_out <= in600;


            when "1001011001" =>
                mux_out <= in601;


            when "1001011010" =>
                mux_out <= in602;


            when "1001011011" =>
                mux_out <= in603;


            when "1001011100" =>
                mux_out <= in604;


            when "1001011101" =>
                mux_out <= in605;


            when "1001011110" =>
                mux_out <= in606;


            when "1001011111" =>
                mux_out <= in607;


            when "1001100000" =>
                mux_out <= in608;


            when "1001100001" =>
                mux_out <= in609;


            when "1001100010" =>
                mux_out <= in610;


            when "1001100011" =>
                mux_out <= in611;


            when "1001100100" =>
                mux_out <= in612;


            when "1001100101" =>
                mux_out <= in613;


            when "1001100110" =>
                mux_out <= in614;


            when "1001100111" =>
                mux_out <= in615;


            when "1001101000" =>
                mux_out <= in616;


            when "1001101001" =>
                mux_out <= in617;


            when "1001101010" =>
                mux_out <= in618;


            when "1001101011" =>
                mux_out <= in619;


            when "1001101100" =>
                mux_out <= in620;


            when "1001101101" =>
                mux_out <= in621;


            when "1001101110" =>
                mux_out <= in622;


            when "1001101111" =>
                mux_out <= in623;


            when "1001110000" =>
                mux_out <= in624;


            when "1001110001" =>
                mux_out <= in625;


            when "1001110010" =>
                mux_out <= in626;


            when "1001110011" =>
                mux_out <= in627;


            when "1001110100" =>
                mux_out <= in628;


            when "1001110101" =>
                mux_out <= in629;


            when "1001110110" =>
                mux_out <= in630;


            when "1001110111" =>
                mux_out <= in631;


            when "1001111000" =>
                mux_out <= in632;


            when "1001111001" =>
                mux_out <= in633;


            when "1001111010" =>
                mux_out <= in634;


            when "1001111011" =>
                mux_out <= in635;


            when "1001111100" =>
                mux_out <= in636;


            when "1001111101" =>
                mux_out <= in637;


            when "1001111110" =>
                mux_out <= in638;


            when "1001111111" =>
                mux_out <= in639;


            when "1010000000" =>
                mux_out <= in640;


            when "1010000001" =>
                mux_out <= in641;


            when "1010000010" =>
                mux_out <= in642;


            when "1010000011" =>
                mux_out <= in643;


            when "1010000100" =>
                mux_out <= in644;


            when "1010000101" =>
                mux_out <= in645;


            when "1010000110" =>
                mux_out <= in646;


            when "1010000111" =>
                mux_out <= in647;


            when "1010001000" =>
                mux_out <= in648;


            when "1010001001" =>
                mux_out <= in649;


            when "1010001010" =>
                mux_out <= in650;


            when "1010001011" =>
                mux_out <= in651;


            when "1010001100" =>
                mux_out <= in652;


            when "1010001101" =>
                mux_out <= in653;


            when "1010001110" =>
                mux_out <= in654;


            when "1010001111" =>
                mux_out <= in655;


            when "1010010000" =>
                mux_out <= in656;


            when "1010010001" =>
                mux_out <= in657;


            when "1010010010" =>
                mux_out <= in658;


            when "1010010011" =>
                mux_out <= in659;


            when "1010010100" =>
                mux_out <= in660;


            when "1010010101" =>
                mux_out <= in661;


            when "1010010110" =>
                mux_out <= in662;


            when "1010010111" =>
                mux_out <= in663;


            when "1010011000" =>
                mux_out <= in664;


            when "1010011001" =>
                mux_out <= in665;


            when "1010011010" =>
                mux_out <= in666;


            when "1010011011" =>
                mux_out <= in667;


            when "1010011100" =>
                mux_out <= in668;


            when "1010011101" =>
                mux_out <= in669;


            when "1010011110" =>
                mux_out <= in670;


            when "1010011111" =>
                mux_out <= in671;


            when "1010100000" =>
                mux_out <= in672;


            when "1010100001" =>
                mux_out <= in673;


            when "1010100010" =>
                mux_out <= in674;


            when "1010100011" =>
                mux_out <= in675;


            when "1010100100" =>
                mux_out <= in676;


            when "1010100101" =>
                mux_out <= in677;


            when "1010100110" =>
                mux_out <= in678;


            when "1010100111" =>
                mux_out <= in679;


            when "1010101000" =>
                mux_out <= in680;


            when "1010101001" =>
                mux_out <= in681;


            when "1010101010" =>
                mux_out <= in682;


            when "1010101011" =>
                mux_out <= in683;


            when "1010101100" =>
                mux_out <= in684;


            when "1010101101" =>
                mux_out <= in685;


            when "1010101110" =>
                mux_out <= in686;


            when "1010101111" =>
                mux_out <= in687;


            when "1010110000" =>
                mux_out <= in688;


            when "1010110001" =>
                mux_out <= in689;


            when "1010110010" =>
                mux_out <= in690;


            when "1010110011" =>
                mux_out <= in691;


            when "1010110100" =>
                mux_out <= in692;


            when "1010110101" =>
                mux_out <= in693;


            when "1010110110" =>
                mux_out <= in694;


            when "1010110111" =>
                mux_out <= in695;


            when "1010111000" =>
                mux_out <= in696;


            when "1010111001" =>
                mux_out <= in697;


            when "1010111010" =>
                mux_out <= in698;


            when "1010111011" =>
                mux_out <= in699;


            when "1010111100" =>
                mux_out <= in700;


            when "1010111101" =>
                mux_out <= in701;


            when "1010111110" =>
                mux_out <= in702;


            when "1010111111" =>
                mux_out <= in703;


            when "1011000000" =>
                mux_out <= in704;


            when "1011000001" =>
                mux_out <= in705;


            when "1011000010" =>
                mux_out <= in706;


            when "1011000011" =>
                mux_out <= in707;


            when "1011000100" =>
                mux_out <= in708;


            when "1011000101" =>
                mux_out <= in709;


            when "1011000110" =>
                mux_out <= in710;


            when "1011000111" =>
                mux_out <= in711;


            when "1011001000" =>
                mux_out <= in712;


            when "1011001001" =>
                mux_out <= in713;


            when "1011001010" =>
                mux_out <= in714;


            when "1011001011" =>
                mux_out <= in715;


            when "1011001100" =>
                mux_out <= in716;


            when "1011001101" =>
                mux_out <= in717;


            when "1011001110" =>
                mux_out <= in718;


            when "1011001111" =>
                mux_out <= in719;


            when "1011010000" =>
                mux_out <= in720;


            when "1011010001" =>
                mux_out <= in721;


            when "1011010010" =>
                mux_out <= in722;


            when "1011010011" =>
                mux_out <= in723;


            when "1011010100" =>
                mux_out <= in724;


            when "1011010101" =>
                mux_out <= in725;


            when "1011010110" =>
                mux_out <= in726;


            when "1011010111" =>
                mux_out <= in727;


            when "1011011000" =>
                mux_out <= in728;


            when "1011011001" =>
                mux_out <= in729;


            when "1011011010" =>
                mux_out <= in730;


            when "1011011011" =>
                mux_out <= in731;


            when "1011011100" =>
                mux_out <= in732;


            when "1011011101" =>
                mux_out <= in733;


            when "1011011110" =>
                mux_out <= in734;


            when "1011011111" =>
                mux_out <= in735;


            when "1011100000" =>
                mux_out <= in736;


            when "1011100001" =>
                mux_out <= in737;


            when "1011100010" =>
                mux_out <= in738;


            when "1011100011" =>
                mux_out <= in739;


            when "1011100100" =>
                mux_out <= in740;


            when "1011100101" =>
                mux_out <= in741;


            when "1011100110" =>
                mux_out <= in742;


            when "1011100111" =>
                mux_out <= in743;


            when "1011101000" =>
                mux_out <= in744;


            when "1011101001" =>
                mux_out <= in745;


            when "1011101010" =>
                mux_out <= in746;


            when "1011101011" =>
                mux_out <= in747;


            when "1011101100" =>
                mux_out <= in748;


            when "1011101101" =>
                mux_out <= in749;


            when "1011101110" =>
                mux_out <= in750;


            when "1011101111" =>
                mux_out <= in751;


            when "1011110000" =>
                mux_out <= in752;


            when "1011110001" =>
                mux_out <= in753;


            when "1011110010" =>
                mux_out <= in754;


            when "1011110011" =>
                mux_out <= in755;


            when "1011110100" =>
                mux_out <= in756;


            when "1011110101" =>
                mux_out <= in757;


            when "1011110110" =>
                mux_out <= in758;


            when "1011110111" =>
                mux_out <= in759;


            when "1011111000" =>
                mux_out <= in760;


            when "1011111001" =>
                mux_out <= in761;


            when "1011111010" =>
                mux_out <= in762;


            when "1011111011" =>
                mux_out <= in763;


            when "1011111100" =>
                mux_out <= in764;


            when "1011111101" =>
                mux_out <= in765;


            when "1011111110" =>
                mux_out <= in766;


            when "1011111111" =>
                mux_out <= in767;


            when "1100000000" =>
                mux_out <= in768;


            when "1100000001" =>
                mux_out <= in769;


            when "1100000010" =>
                mux_out <= in770;


            when "1100000011" =>
                mux_out <= in771;


            when "1100000100" =>
                mux_out <= in772;


            when "1100000101" =>
                mux_out <= in773;


            when "1100000110" =>
                mux_out <= in774;


            when "1100000111" =>
                mux_out <= in775;


            when "1100001000" =>
                mux_out <= in776;


            when "1100001001" =>
                mux_out <= in777;


            when "1100001010" =>
                mux_out <= in778;


            when "1100001011" =>
                mux_out <= in779;


            when "1100001100" =>
                mux_out <= in780;


            when "1100001101" =>
                mux_out <= in781;


            when "1100001110" =>
                mux_out <= in782;


            when "1100001111" =>
                mux_out <= in783;


            when "1100010000" =>
                mux_out <= in784;


            when "1100010001" =>
                mux_out <= in785;


            when "1100010010" =>
                mux_out <= in786;


            when "1100010011" =>
                mux_out <= in787;


            when "1100010100" =>
                mux_out <= in788;


            when "1100010101" =>
                mux_out <= in789;


            when "1100010110" =>
                mux_out <= in790;


            when "1100010111" =>
                mux_out <= in791;


            when "1100011000" =>
                mux_out <= in792;


            when "1100011001" =>
                mux_out <= in793;


            when "1100011010" =>
                mux_out <= in794;


            when "1100011011" =>
                mux_out <= in795;


            when "1100011100" =>
                mux_out <= in796;


            when "1100011101" =>
                mux_out <= in797;


            when "1100011110" =>
                mux_out <= in798;


            when "1100011111" =>
                mux_out <= in799;


            when "1100100000" =>
                mux_out <= in800;


            when "1100100001" =>
                mux_out <= in801;


            when "1100100010" =>
                mux_out <= in802;


            when "1100100011" =>
                mux_out <= in803;


            when "1100100100" =>
                mux_out <= in804;


            when "1100100101" =>
                mux_out <= in805;


            when "1100100110" =>
                mux_out <= in806;


            when "1100100111" =>
                mux_out <= in807;


            when "1100101000" =>
                mux_out <= in808;


            when "1100101001" =>
                mux_out <= in809;


            when "1100101010" =>
                mux_out <= in810;


            when "1100101011" =>
                mux_out <= in811;


            when "1100101100" =>
                mux_out <= in812;


            when "1100101101" =>
                mux_out <= in813;


            when "1100101110" =>
                mux_out <= in814;


            when "1100101111" =>
                mux_out <= in815;


            when "1100110000" =>
                mux_out <= in816;


            when "1100110001" =>
                mux_out <= in817;


            when "1100110010" =>
                mux_out <= in818;


            when "1100110011" =>
                mux_out <= in819;


            when "1100110100" =>
                mux_out <= in820;


            when "1100110101" =>
                mux_out <= in821;


            when "1100110110" =>
                mux_out <= in822;


            when "1100110111" =>
                mux_out <= in823;


            when "1100111000" =>
                mux_out <= in824;


            when "1100111001" =>
                mux_out <= in825;


            when "1100111010" =>
                mux_out <= in826;


            when "1100111011" =>
                mux_out <= in827;


            when "1100111100" =>
                mux_out <= in828;


            when "1100111101" =>
                mux_out <= in829;


            when "1100111110" =>
                mux_out <= in830;


            when "1100111111" =>
                mux_out <= in831;


            when "1101000000" =>
                mux_out <= in832;


            when "1101000001" =>
                mux_out <= in833;


            when "1101000010" =>
                mux_out <= in834;


            when "1101000011" =>
                mux_out <= in835;


            when "1101000100" =>
                mux_out <= in836;


            when "1101000101" =>
                mux_out <= in837;


            when "1101000110" =>
                mux_out <= in838;


            when "1101000111" =>
                mux_out <= in839;


            when "1101001000" =>
                mux_out <= in840;


            when "1101001001" =>
                mux_out <= in841;


            when "1101001010" =>
                mux_out <= in842;


            when "1101001011" =>
                mux_out <= in843;


            when "1101001100" =>
                mux_out <= in844;


            when "1101001101" =>
                mux_out <= in845;


            when "1101001110" =>
                mux_out <= in846;


            when "1101001111" =>
                mux_out <= in847;


            when "1101010000" =>
                mux_out <= in848;


            when "1101010001" =>
                mux_out <= in849;


            when "1101010010" =>
                mux_out <= in850;


            when "1101010011" =>
                mux_out <= in851;


            when "1101010100" =>
                mux_out <= in852;


            when "1101010101" =>
                mux_out <= in853;


            when "1101010110" =>
                mux_out <= in854;


            when "1101010111" =>
                mux_out <= in855;


            when "1101011000" =>
                mux_out <= in856;


            when "1101011001" =>
                mux_out <= in857;


            when "1101011010" =>
                mux_out <= in858;


            when "1101011011" =>
                mux_out <= in859;


            when "1101011100" =>
                mux_out <= in860;


            when "1101011101" =>
                mux_out <= in861;


            when "1101011110" =>
                mux_out <= in862;


            when "1101011111" =>
                mux_out <= in863;


            when "1101100000" =>
                mux_out <= in864;


            when "1101100001" =>
                mux_out <= in865;


            when "1101100010" =>
                mux_out <= in866;


            when "1101100011" =>
                mux_out <= in867;


            when "1101100100" =>
                mux_out <= in868;


            when "1101100101" =>
                mux_out <= in869;


            when "1101100110" =>
                mux_out <= in870;


            when "1101100111" =>
                mux_out <= in871;


            when "1101101000" =>
                mux_out <= in872;


            when "1101101001" =>
                mux_out <= in873;


            when "1101101010" =>
                mux_out <= in874;


            when "1101101011" =>
                mux_out <= in875;


            when "1101101100" =>
                mux_out <= in876;


            when "1101101101" =>
                mux_out <= in877;


            when "1101101110" =>
                mux_out <= in878;


            when "1101101111" =>
                mux_out <= in879;


            when "1101110000" =>
                mux_out <= in880;


            when "1101110001" =>
                mux_out <= in881;


            when "1101110010" =>
                mux_out <= in882;


            when "1101110011" =>
                mux_out <= in883;


            when "1101110100" =>
                mux_out <= in884;


            when "1101110101" =>
                mux_out <= in885;


            when "1101110110" =>
                mux_out <= in886;


            when "1101110111" =>
                mux_out <= in887;


            when "1101111000" =>
                mux_out <= in888;


            when "1101111001" =>
                mux_out <= in889;


            when "1101111010" =>
                mux_out <= in890;


            when "1101111011" =>
                mux_out <= in891;


            when "1101111100" =>
                mux_out <= in892;


            when "1101111101" =>
                mux_out <= in893;


            when "1101111110" =>
                mux_out <= in894;


            when "1101111111" =>
                mux_out <= in895;


            when "1110000000" =>
                mux_out <= in896;


            when "1110000001" =>
                mux_out <= in897;


            when "1110000010" =>
                mux_out <= in898;


            when "1110000011" =>
                mux_out <= in899;


            when "1110000100" =>
                mux_out <= in900;


            when "1110000101" =>
                mux_out <= in901;


            when "1110000110" =>
                mux_out <= in902;


            when "1110000111" =>
                mux_out <= in903;


            when "1110001000" =>
                mux_out <= in904;


            when "1110001001" =>
                mux_out <= in905;


            when "1110001010" =>
                mux_out <= in906;


            when "1110001011" =>
                mux_out <= in907;


            when "1110001100" =>
                mux_out <= in908;


            when "1110001101" =>
                mux_out <= in909;


            when "1110001110" =>
                mux_out <= in910;


            when "1110001111" =>
                mux_out <= in911;


            when "1110010000" =>
                mux_out <= in912;


            when "1110010001" =>
                mux_out <= in913;


            when "1110010010" =>
                mux_out <= in914;


            when "1110010011" =>
                mux_out <= in915;


            when "1110010100" =>
                mux_out <= in916;


            when "1110010101" =>
                mux_out <= in917;


            when "1110010110" =>
                mux_out <= in918;


            when "1110010111" =>
                mux_out <= in919;


            when "1110011000" =>
                mux_out <= in920;


            when "1110011001" =>
                mux_out <= in921;


            when "1110011010" =>
                mux_out <= in922;


            when "1110011011" =>
                mux_out <= in923;


            when "1110011100" =>
                mux_out <= in924;


            when "1110011101" =>
                mux_out <= in925;


            when "1110011110" =>
                mux_out <= in926;


            when "1110011111" =>
                mux_out <= in927;


            when "1110100000" =>
                mux_out <= in928;


            when "1110100001" =>
                mux_out <= in929;


            when "1110100010" =>
                mux_out <= in930;


            when "1110100011" =>
                mux_out <= in931;


            when "1110100100" =>
                mux_out <= in932;


            when "1110100101" =>
                mux_out <= in933;


            when "1110100110" =>
                mux_out <= in934;


            when "1110100111" =>
                mux_out <= in935;


            when "1110101000" =>
                mux_out <= in936;


            when "1110101001" =>
                mux_out <= in937;


            when "1110101010" =>
                mux_out <= in938;


            when "1110101011" =>
                mux_out <= in939;


            when "1110101100" =>
                mux_out <= in940;


            when "1110101101" =>
                mux_out <= in941;


            when "1110101110" =>
                mux_out <= in942;


            when "1110101111" =>
                mux_out <= in943;


            when "1110110000" =>
                mux_out <= in944;


            when "1110110001" =>
                mux_out <= in945;


            when "1110110010" =>
                mux_out <= in946;


            when "1110110011" =>
                mux_out <= in947;


            when "1110110100" =>
                mux_out <= in948;


            when "1110110101" =>
                mux_out <= in949;


            when "1110110110" =>
                mux_out <= in950;


            when "1110110111" =>
                mux_out <= in951;


            when "1110111000" =>
                mux_out <= in952;


            when "1110111001" =>
                mux_out <= in953;


            when "1110111010" =>
                mux_out <= in954;


            when "1110111011" =>
                mux_out <= in955;


            when "1110111100" =>
                mux_out <= in956;


            when "1110111101" =>
                mux_out <= in957;


            when "1110111110" =>
                mux_out <= in958;


            when "1110111111" =>
                mux_out <= in959;


            when "1111000000" =>
                mux_out <= in960;


            when "1111000001" =>
                mux_out <= in961;


            when "1111000010" =>
                mux_out <= in962;


            when "1111000011" =>
                mux_out <= in963;


            when "1111000100" =>
                mux_out <= in964;


            when "1111000101" =>
                mux_out <= in965;


            when "1111000110" =>
                mux_out <= in966;


            when "1111000111" =>
                mux_out <= in967;


            when "1111001000" =>
                mux_out <= in968;


            when "1111001001" =>
                mux_out <= in969;


            when "1111001010" =>
                mux_out <= in970;


            when "1111001011" =>
                mux_out <= in971;


            when "1111001100" =>
                mux_out <= in972;


            when "1111001101" =>
                mux_out <= in973;


            when "1111001110" =>
                mux_out <= in974;


            when "1111001111" =>
                mux_out <= in975;


            when "1111010000" =>
                mux_out <= in976;


            when "1111010001" =>
                mux_out <= in977;


            when "1111010010" =>
                mux_out <= in978;


            when "1111010011" =>
                mux_out <= in979;


            when "1111010100" =>
                mux_out <= in980;


            when "1111010101" =>
                mux_out <= in981;


            when "1111010110" =>
                mux_out <= in982;


            when "1111010111" =>
                mux_out <= in983;


            when "1111011000" =>
                mux_out <= in984;


            when "1111011001" =>
                mux_out <= in985;


            when "1111011010" =>
                mux_out <= in986;


            when "1111011011" =>
                mux_out <= in987;


            when "1111011100" =>
                mux_out <= in988;


            when "1111011101" =>
                mux_out <= in989;


            when "1111011110" =>
                mux_out <= in990;


            when "1111011111" =>
                mux_out <= in991;


            when "1111100000" =>
                mux_out <= in992;


            when "1111100001" =>
                mux_out <= in993;


            when "1111100010" =>
                mux_out <= in994;


            when "1111100011" =>
                mux_out <= in995;


            when "1111100100" =>
                mux_out <= in996;


            when "1111100101" =>
                mux_out <= in997;


            when "1111100110" =>
                mux_out <= in998;


            when "1111100111" =>
                mux_out <= in999;


            when "1111101000" =>
                mux_out <= in1000;


            when "1111101001" =>
                mux_out <= in1001;


            when "1111101010" =>
                mux_out <= in1002;


            when "1111101011" =>
                mux_out <= in1003;


            when "1111101100" =>
                mux_out <= in1004;


            when "1111101101" =>
                mux_out <= in1005;


            when "1111101110" =>
                mux_out <= in1006;


            when "1111101111" =>
                mux_out <= in1007;


            when "1111110000" =>
                mux_out <= in1008;


            when "1111110001" =>
                mux_out <= in1009;


            when "1111110010" =>
                mux_out <= in1010;


            when "1111110011" =>
                mux_out <= in1011;


            when "1111110100" =>
                mux_out <= in1012;


            when "1111110101" =>
                mux_out <= in1013;


            when "1111110110" =>
                mux_out <= in1014;


            when "1111110111" =>
                mux_out <= in1015;


            when "1111111000" =>
                mux_out <= in1016;


            when "1111111001" =>
                mux_out <= in1017;


            when "1111111010" =>
                mux_out <= in1018;


            when "1111111011" =>
                mux_out <= in1019;


            when "1111111100" =>
                mux_out <= in1020;


            when "1111111101" =>
                mux_out <= in1021;


            when "1111111110" =>
                mux_out <= in1022;


            when others =>
                mux_out <= in1023;


        end case;

    end process selection;


end architecture behavior;


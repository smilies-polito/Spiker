library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_784x128_exc_ip is
	port(
		clka	: in std_logic;
		addra	: in std_logic_vector(9 downto 0);
		douta	: out std_logic_vector(511 downto 0)
	);
end entity rom_784x128_exc_ip; 

architecture behavior of rom_784x128_exc_ip is

	type rom_type is array(0 to 784) of std_logic_vector(511 downto 0);

	constant mem	: rom_type := (
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00001111000111100001111000010000000011100000111100001110111100000000000000000000000111110001000011110000000000000001111000000000000100001111000011110000000100001110000100000000111111110001000000010000001000011111111100101111000000000000000000000000000000000000000011110000111100011110001000000001000011100001000000000001000100010000000111110000111100000000000100010000000100000000000000010000111111110000000000000010000100010000000000001111000000001111000000000000111000001111111100010001000100001111000100011111",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000011110000111100000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000",
		"00000000000000001111000000000000000000001111111100000000111100010000000000000000000000001111000100010000000100000001000000000000000000000001000000000000000000000000000000000000000000010000111100000000111111111111000100000000000000000000000011110000000000010000000100000000000000000000111100000001000000001111000000001111000000011111000011110001000000000000000100011111111100000000111100000000000000010000000000000001000000010000000000010000111100000001111100000001000000010000000000000000000000000000000100000001",
		"00000000000011110000111100000000000011110000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001111000000000000000000000001000000000000",
		"00000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000",
		"00000000000000000000000000000000000000100000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000100000000000000001000000000000000000001111000000000000000000000000000000010000000000000000000011110001000100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011110000000100000000000000000000111100000000111100000001000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000100010000000100000001000000000000",
		"00000000000000000000000011110000000000000000000000010001000000001111000000000000000000000000000000000000000000000000000000000000000011110001000100001111000000000000000000001111000000000000000000000000000011110000000000001111000000000000000000000000000000010000000000000000111100000000111100010001000000000000000100000000000000000000000000000000000111110000000100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000010000000000000000000111110000",
		"00000000000000000000000000000000000000010000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000011110000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
		"00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000010000000011110000111100010000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000001000000000001000000000000000000010000000000010000000011110000111100000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000010001111100001111000000010000111000100000000000001111000000011110000000001111000000010000000000000000000000000000000100001111000000000000000100000000000000000000111100000000000000000000000100000000000000001111111100001111000011110001000100010000111100000000000000000000000000010010000000000001000000000001000000000000000011111111000000000000000100001111000000000000111100010000000000000001000000000000000000000000000000000000000000000010000000000000111100001111000000000000000000000000000000000000",
		"00000000000000000001111100000000000011111111111000010001111100100000000000011111001000001110000000000000000000000000111100000000000111110000000000000000001000000000000000000000111111110000000000000010000100000000000000000000111100001111111100000010000000011110000000000000000000010000000000010010000000000001000000000001000000000001111111111111111111110001000100000000000000000000111100010000000011110001111100000000000000011111000011111111111100000001000000000000000011111111000000011111000000010000000100000000",
		"00000000000000000000111100000000000000000000111100010001111100010000000000001111000100001111000000000000000000000000111100000000000011110000000000001111000100000000000000000000111111110000000000010001000111100001000000000000111100000000000000000001000000011111000000001111111100000000000000010010000000000000000000010000000000000001111111111111111111110001000100000000000000010000000000010000000000000000111100000000000000011111000000001111000000000010000000000001000011110000000000011110000000000001000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000",
		"00000000000000000000111100000000000000011111000000000001000000010000000000000000000000001111000000000000000000000001000000000000000000000000000000000000000000000000000000000000111100000000111100010000000011110000000100000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000111110000000100001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000",
		"00001111000100001111111111110000000000100000000000000001000000011111000011110000000000000000000100000001000100000001000000010000000011110001000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000100000000000100010000000000001111000000001111111100000001000000001111000100000000000000000000000000000000000011110001000100000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000100011111000000000000000011110001",
		"00000000000000001111000011110000000000010000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000011110001000000000000000000000000000000000000000000000000000000000000111100000001000000000000000000001111000100000000000000000000000000001111000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000001111000000000000000011110001",
		"00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000111111110000000000000000111100000000000000000000000000000000000000000000000011110000000100000000000000000000000000000000000000000000000100000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011110000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000001111000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000111000010001000100010000000000010001000000001111111100000000000000000000000100000001001000010001111100000000111111110000111100001111111100010000111100001111111100010000111100010000000111110000000100000000000100000000000000000000000000010000000100011111111111111111000000000001000000001111000000000000000100011111000000000000000011110000000100011111111100000001111100010001000100010000000100000001111100010001111100001111111111110001111100010001111100001111000100011111000100000000000111110001",
		"00000000000000000000111100000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000010000000000000000000000100000000000000000000000000000000000001111000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000011110000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000001111000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000001111000000000001000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000100000000111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000111100000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001111000000001111000000000001000000000000",
		"00000000000000000000000000000000000000000000111100000000000000001111000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000011111000000000000000000000000000100000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000010000000000000000000000000000",
		"00001111000111100000000000000000000000000000111100000000000000000000000000000000001000000000000011110000000000000000000000000000000000000000111100001111000000000000000000010000111100000000000100010000000100001110000000011111000000010001000000000000000000000000000100001111000000000000000100000000000011110000000000000000000000010000000100000000111100000000000000001111000000000000000000000000000000000000000000010000000000010000000000001111000000000000000100010000000000000000000000000000000000010000000000011111",
		"00000000000011110000000000000000000100000000111100000000000000010000000011110000000100001111111111110000000000000001111100000000000000000000111100000000000000000000000000010000111100001111000000010000000100011111000000001111000000000000000000000000000000010000000000000000000000001111000100000000000000000000000000000000000000010000000011110000111111100000000000000000000000010000000000010001111100000000111100010000000000100000000100000000000000000001001000000001111100000000000000000001000000100000000000000000",
		"00010001000000001111111100000000000100000000111000010000000000000000000011110000000100001111000011110000000000010001111100000001000011100000000000001111000000000000000100001111111100001111000000000000000000000000000111100000000100000000000000000000000000010000000100000000111000001111000111110000000000000000000100000001000000011111111111100000000011110000000100010000000000010000000000100000000000000000000000000001000000010000000111111111111100000000000100000001111100001110000000010000000000011111000000000000",
		"00001111000011110000111000010000000100000000111000000000000000000000000000000000000000011111000011110000000100010000000000000001000011100000000000000000111100100000000000000000000000001111000000010000000000010000000000000000000100000001000000000000000100000000000100000000000000001111000000000000000000010001000000000010000100001111000011110000000111110000001000000000000000000001000100000001000000001111111100000001000000010000001000001111000000000000000100010001000000001110000000100000000000000000000100010000",
		"00001110001000000000000000100000000011110001000000000000111100001111000000000000111100010000000100001111001000000000000100000010000111100000000000000000111000100001000000101110000000001111000000001111000000010000000000000000000000010001000011111111001000000000000000000000000000001111000000011111000000000010000000000010000000000000000000000000001000000000001000001111000000010001000000000000000100000000000000010000000000000001001000000000000111110001000100000000000000011101000000000000000000001111000100000000",
		"00001110000100000000000000010000000011110000000000000000000000001111000000000010000000001111000100001111001000000001000000000010000011010000000000000000111100010001000100101111000000011111000000001110000000011111000000000000000000000000000011111111000100000000000000000000000000001111000000000001000000000000000011110001000000011111000100000000000100000000000100000000000000100000000100000000000100001111000000010000000000100000000000011111000000000000000000010001000000011111000100000000000100001111000000000000",
		"00010000000000001111111100010000000111110000000100010000000000011111000011110001000000000000000000010000000100000001000000000000000000000000000000000000111100000010000100000000000000000000000000011110000000010000000000000000000011110000000000001111000100000000000000000000000000001111000000000001000000001111000111110010111100000000000100000000000000001111000100010000111100010001000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000001111000011110000000000011110000000010000",
		"00000000000000001111000000100000000111110000000000100000111100011111000011110000000000000000000000010000000100000001000000000000111100000000000100000000000000000010000000001111111100000001111100001110000000100000000000000000000000000000000000000000000100001111000000000000000000000000000000000001000000001111000000000010111100000000000100000000000000000000000000010000000000000001111100000000000000000000111100000000000000010001000011110000000000000001000000000000000000000000000000000000000000011110000100000000",
		"00001111000000010000000000010000000100000000000100000000000000001111000011110000000000000000000000010000000000000001000000000010111100000001000000000000000000000000000000000000111100000001000000001110000000010001000000000000000100000000000000001111000000001111111100001111000000000000000000000000000011111111001000000001111100000000000100000000000000010000000000000000111100010000000000001111000000000000000000000000000000010001000000000000000000000000000000001111000000000000000111111110000000010000000000000001",
		"00001110000000011111111100000000001000001111000000000000000000001111000011110000000000000001000000010000000000000010000000000001000011110000000000000000000000000001000000000001000000000001111100001111000111110000000100000000000111110001000000001111000000001111111111111110000000001111000000000000000011100000000000000001111100001111000000000001000000000000000000000000000000010000000000000000000000010000000000000000000000010000111100010000000000000000000100000000000000001111000100011101000000000001000000000001",
		"00000000000100011111111100000000000000011101000000010000000000001110000000000000111100010000000000000001000100010001000000000001000000000001111100000000000000000010000000000000111100000001111000001110000000000001000000010000000000001111000000001111000000000000000000001111000000000000000000000000111111111111000011111111111100000000000000000000000000010000000100001111111100000000000000000000000000010000001000011111000000100000111100000000111100000000000000000000000000001111000100011110000000000010000000000001",
		"00001111000000001111111100000000000000011111000000010001000000001111000011110000111100000000000000000001000000000001000000000000000011110001000000000000000000000010000000001111111100000000111000000000000000000000000000010000000000000000000000001111000100000001000000000000000000000000000000000000111100001110000011100000000000010000000011110000000000000000000100000000111100010000000000000000000000000000000100000000000000010000000000000000000000000000000000000000111100001111000000011111000000000000000000000000",
		"00000000000011110000111100000000000000000000000000010001000000010000000011110000000000000001000100000001000100000000000100000000111100000000000000000000000000000000000000001111000000000000111100001111000011110000000000000000000000000000000100000000000100010001000100000000000000000000000000010001000000001110000100001111000000001111000000000000000011110000000100000000111100000000000000010000000000010000000100000000000000010000000000001111000000000000000000000000111100001111000000101110000000000000001011110001",
		"00000000000000001111000000000000000000000000000000000001000000001111000011110000111100000000000000000001000100000000000000010000000000000000000000000000000000000000000000000000111100000000000000000000000011110000000000011111000000001111000000000000000000000000000000000000000000000000000000000000000000001111000100000000000000000000000000000000000000000000000000000000111100000000000000010000000000000000000000000000111100000000000000010000000000000001000000000000000000010000000000011111000000000000000111110001",
		"00000000000000000000111100000000000000001111000000000000000000010000000011110000000000000000000000000000000100000001000000010000111111110000000000001111000000000000000000000000000000000000000000000000000000001111000100000000000000000000000000000000000000010000000000001111000000000000000000000000000000000000000100000000000000010000000100000000000011110000000000000000000000000000000000000000000000000000000000000000000000010000000000011111000000000001000000000000000000001111000000010000000000001111000000000000",
		"00000000000000000000000000000000000000000000111100000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001111000000010000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000111100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"11111111000000010000001000011111000100011111111111110000000111111111000111110000111100000001000000100000000100000001000100000001000100011110000011110001000011100001000000001111000000000000000100010000111100100001000000000001111000010001000100000010000011110001000000010001000011110010000000001111000000010000111100000001000000100001111100000000111000010001001000101111000000000010000000011111111000000000000000001111000100000001001000000001000100010010000111111111111100101110111111110001000000010000000011111111",
		"00001111000000000000000000010000000000010000000000000000000000001111000011111111000000000000111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000111100000000111100010000000000000000111100000000000000000000000000000000000000000000000000000000000000010000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000011111111",
		"00010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000000000000000000000000000000000111100000000000000000000000000000000000000001111000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100011111000000000000000000000000000000000000111100000000000000000000000000010000000100010000000000000000000100000000111100000000000000000000000000000000000000000000000000000000000000000001",
		"00000000000000000000111000000000000111110000000000000000111100000000000000000000000000000000000111110000000100000010000000000000111100000000000000000000000000000000000100000000111100001111000000010000000100000000000100001111000100000000000000000000000100001111000000000000111100001111000011110001000000000000000111110000000000000000000011110000000011111111000000010000000000001111000000010001000000000000000000010000000000010000000000000000000011110001000000000000000000000000000000000000000000010000000000000000",
		"00010000000000001111111000010000000111110000000000100000111100010000000011110000000000000000000100000000000100000010000000000000111111110000000000000000000000000000000000000000000000000000000000010000000100000000000100011110000100000000000000000000000000000000000000000000111100001111000000000001000000000000000000000000000000011111000011110000111100000000000100010000000100010000111100000000000000000000000000000000000000010000000100000000000000000000000100000000111100010000000100000000000000010000000000000000",
		"00010000000000000000111000100000000000000000111100100000000000000000000011110000000011111111000011110000001000010010000000000000111011100000000100000000000000010000000100001111000000000000000000000000000000000000000000011111000100000000000000000000000100000000000000001111111100000000000011110010000000001111001000000000000000000000000000000000000011110000001000001111000000001111111100000001000000001111000000100000000000000000000100000000000000000000000011110000111100010000000100000000000000000000000011110000",
		"00000000111100000000110100000000000011110000000000010000111100100000000000000000000011111111111100000000000000000010111100000000110111110000000000000001000000011110001011111111111100000000000000000000111100000010000000100000000000000000000000000000000000010000000011111110111100000000000011110011111100001110001000000000000000010000000000001111000011101111001100010000000000011110111100010001000000000000000000100010000000000000000000000000000011110010001011110001111100001111000000000001000000011111000000011111",
		"00000000111100000000111100000000000000000000111100000000000000010000000100000001000011110000000000000000111100000000111100001110111111100000000000000000000000001111000000000000110100000000000000000000000000000000000000111110000100000000000000000001000000100000000011111111111100010000000000000000000011110000000100000000000000010000000000001110111111010000000000000001000000100000111100100000111100000000000000000001000000010000000000100000000000000010001000010000111000001110000100000000000100011111000100011111",
		"00000000111000000000000000001111000000010000000000000000000100010000000000000001111000000000000011111111000000000000111111111111111111100001111100000001000000001111000000010001111100000000000000000000000000000000000000101111000100000000111100010000000000011111000011111111000000000000000000000000000000000000001000000000000000000000000011110000111111101111111100000001000000011110111100011111000000010000111100000000000000010000000000100000000000000001000100100000000011111111000011110000000000000000000100001111",
		"00010000111111110000111100000000000000000000111000010000000000000001000000000001111000000000111100000000000000000000111111110000111011110001000000000000000000000000000011110000000000000000000000000000000000000000000000011111000100000000111100010000000000011110000011100000000000000000111100000000111000000000001100000001000000000000000000001110000011111111000000010000000000001101000000011111000000000000111000010001000000001111000000010000000000000000000100010010000011111110000000000000000100000000000000000000",
		"00010000111100000000000000001111000111110000000000010000000000010000000000000001000000001110111100001111000000010000000000000000111111110010111100000000000000010001000000000000000011110001000000010001111100010000000000011110000000010000111100011110000000101111000011111111000000000001000000000000111000000001001000000001000000010000000000001110000011111111000000010001000000011110000000011111000000000000111100100000000000001111000100010000000000000001001011110001111000001110000000000001000000010000000000011111",
		"00000000111100001111111100000000000111100000000100000000111100011111000111110001000000011100000000010000000000010000000100010001000011010001000000000000000000100001000100000000111100000000000000000000111100000000000000011111000000000000111100001101000000011111000000001111000000001111111100000000111100000000000011100000000000000000001000000000000100000000001000000000111100101111000000001111000000000001000000100000000000010000000000010000000000000000000100000000110100000000000011110000000100010000000000000000",
		"00000001111100000000000000000000000011010001000100000000111000000000000000000000000000010000000100010000000000000000000100000000000011010001001000000000111100010001001000000000000000000000000000010000111100000000000000100000000000000001000000001101000000011100000000000001000000001111000000000001111100000000000111110000111100001111000000000000000000001111000100000000000000000000111100000000000100000000000000100000000000000000000000000000000000000000001000000001111100000000000000001111000000000000000000010000",
		"00000000000000000000000000000000000111010000000000010000111100010000000000000000000000100000000000000000000000000001000100001111000011110000000100000000000000000001001000000000000000000000000000000000111100010000000000100000000000000001000000001110000000001100000100000001000000010000111111110000111100001110000011010000111000000000000100000000000000001110000000000000000000000000111100000000000100000000111100100000000000000000000111110000000000000000000000000000000000000000000100000000000000001111000000001111",
		"00000000000100000000000000010000001011110000000100100000000000010000000000000000000000010010000000000000111100000000000000001111000011110000000000000000000000010001000100000000111100001111000000000000111100000000000000000001111111110001000000001110000000001101000111110001000000010000111111110001000000001111000011100001111100000000000111110000000011111111000100000000000000000000111100000000000100000000000000010000000000000000000000001111000000000000000100000000000000010000000000000000000000001111000000010000",
		"00000000000000000000000000010000001000011111000000010000111000000000000000000000000000010001111100000000000000000000000000000001000000000001000000000000000000010010000100000000111100000000000000000000111100000000000000000010000000000001000000001111000000001110000011110001000000010000000000000000000000011111000100000000000000000000000000000000000000010000000000000000111100010001000000001111000000000000000000000000000000000000000011110000000011110000000000000000000000010000000100001110000000000000000000010000",
		"00000000000000001111000000011111001100010000000100000000000000101111000000000000000000001111111100000000111100000000111100010011000000100001000000000000000000010010000000000000111100000000000000000000111000000001000000000001000000010001000000001110000011111111000011110000000000000000000000001111000000001111000100001111000000000000000000000001000000010000000000000000111000000000000100001111000000000000000000011111000100000001111100000000000011100000000000000000000000000000000100001101000000000010000100000000",
		"11110001000100001111000000001110000100011110000100000000000100000000000000000000000000010000000000000000111111110001111000100010000000000000111000000000000000000010000000000000000000010000000011110000111100010001000100000000000000100000000000001110000000000000000011110001000000000000000000001101111100001101000000010000000000000000000000000000000000100000000000001111111100010000000000010000000100000000000000001111001000000000000011110000000111110000000000010000111100000000001000011110000000000000000000000001",
		"11110011000000000000000000001111111100011111000100010001000000010000000000000000111100010001000000000000000011110000000000000001111011110000000000000000000000000011000000000000000000010001000011110000111000000010000100000000000000010000000000001111000000000000111111110001000000000000000011110000111100010000000000000000000100000000000000000000000000101111111100000000111100011111000100010000000100000000111100000000000111110000000000000000000000000010000100010000000000000001001000001110000000000000000000100000",
		"00000000000000000000000100001111000000000001000000010000111100010000000000000000000000010001000000000000000000000001000000000001000011110000000000000000000000010001000000000000000000010001000000000000111111110000000000000000000100000000000000010000000000010000000000001111000000000000000000000001000000001110000000000000000000000000000100000001000000010000000000000000111100010000001000010000000000010000000100000001000100000000111100010000000000000000000000000000111111110001001000001110000000001111000100000001",
		"00001111111100000000001000000000000100000000000000000000000000000000000011110000000100000001000000000001000000000000000000000001000011111111000100000000000000010010111100001111000000100000000000001111000011110001000000000000000000000000000000001111000000000000000000000000111100000000000000010000000000000000111111110000111000000000000111100010000000100000000000000000111100010000000100000000000000100000000100000000000000000000000000010000111100000000000000000000111100000000000100001111000000001111000000000001",
		"00011111000000000000000111110000000100000000111100000001000000010000111100000000000100000000000000000010000000100001000100000000000011110000000000000000000000000001000000000000000000010000000000001110000000000001000011111111000100000000000000000000000000100000000000001111000000000000000000000000000000001111000000000000111000011111000011110001000000000001000000000000000000000001000000000000000000100000000100010000111000000000000000000000000000000001000000010001111100000000000000000000000000000000000011110001",
		"00010000000000000000000000001111000100000000000000000000111100000000000000000000001000001111000000000010000000000001000000000000000000000000111100000000000000000000000100001111000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111000000000000000000101111000011100000000000000000000000000000000000000000000000000000000000000000000100000000111100000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001111111100000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000100001111000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000001000000000000000000000000111100010000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000010000111100000001000000000000000000000000000000001110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000111100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000111100011111000000000000111000000001000000000000000000000001000011111111000000000001000100000000000100000001000000000000000000010001000011110000000000000000000000000000000000000000111100000001000000010001000000000000000000000000000011110000000011110000000000000000000000000001000000001111000000000000000000010000000011110000000011110000000111110000000000001111000000000000000000000000000000000000000011110000000000001111000100000001000000000000000000000000000000000000000000010000111111111111",
		"11111111000100000000001000011110000100010000000011100000000100001111000100000000000000000001000000001111000100000010000100000001000100101111000011110001000011110001111100001110000000000000000100010000000000100001000000000000111100010001000111110010000011100001000000100001000011110001000000001111000000000000111100010000000000100001111000001111111000010010001000011111111111110001000000011111111100000000000000000000000000000001000100000001001000100010000011101111000000011111111111110010000000010000000011101111",
		"11110000000000011111000000011111000000000000000000000000000100000001000000000000000000000000111100000000001000000000000000000001000000000001000000000001000011110001000000001111000000000000000011110000111100010010000000010000111100010000000000000000000011110000111100000000000011110001000000000000000000000000000000010000000000010001000000000000111100000001000000000000000011110001000000010000111100000000000000010000111100000000000100000000000100010001000100000000000000000000111100000010111100000000000011111111",
		"00010000000000000000000000000000000000001111000000010000000000010000000000000000000000001111000100010001000100000000000000000001000000000001000000000000111100000001000000000000111100001111111100000000111100000000000100010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000011110000000000000000000000000000000000000000000000010000000000010000111100000000000000000000000000000001000000000001000000010000111100000000000000000000111100000000",
		"00010000000000000000000000000001000000000000000000000000000000000001000000000001111100001111000100000000000100000001000000000000111011110000000000001111111100000001000100000000000000001111111100010000000100000000000000010001000100000001000100000000000100001111000100010000111100001111000011110000000000001111000000010000000000010000000000001111000011111111111100010000000100001111111100100000000000011111111100000000000000000000000000001111000000000000000100000000000000010000111100000000000100010000000000000000",
		"00000000000000000000000000010000000000000001000000000000000000000001000000000001111111111110000000001111000000000001000000000000110111110000000000000000111000000000000100000000000000010000000000000000000100001111000000000000000100010010000100000000000100000000000000000000000000000000000000000000000000001111000000010000000000010000111100001111000000000000000000010000001000000000000000010000111100000000111100000000000000000000000100000000000000000000001000000000000000000000000000000000000100000000000000001111",
		"00000001111111110000111100000000000000010000000000000000000000010010000100000010000011100000111111110000000000010000111100001111111000000000111100000000000000000000000000000000000000100000000000000000000000000000000000000001000100000001000100000001000100000000000000000000000000100000111100000001000000000000000011110000000000010000000000011110000000000000000000010000001100000000000000000000111100000000111100000000000000001111000000011110000000000000001011110000000000000000000011110001000100000000111011111111",
		"00000000111100000000000000001111000100100000000000001111111000000000000111100001111111100000000000000000000000000001111100001111111100000000110100000000000000000000000000000000111000010000000000100001000000000000000100010000001000000001000100000000000000010000000000000000000000011111000011110000000000001110000111010000000000010000111100000000000111111111001000010000000100011111000000000000111100000001000000000000000000011111111100011110000000000000000000000000000000000000111111110001001000000000000011111111",
		"00000000111100001111000000001110000100010000000000001111110100010000000100000001111000000000000000001111000000000000000000001111111111100001111000000000000000010000000000010001111100010000000000000001000000000000000100001111000100000001000000000000000000010000000000000000000000001110000000000000111100001110000011010000000000010000000000000000000100001111000000010000000000011111000000001111000000010001000100000000000000011111000000000000111100000001000000000000000000000000000000000000001000000000000000000000",
		"00000000111100000000000000001110000100010000000000011110111000010000000111110011111111110000000000001111000100000001000000000000111111100001110100000000000000000000000000000000111100010000000000010001000000010000000000000000000111110000000000000000000000010000000000000001000000001111000011100000111000001110000111010000000000010001000000000000000000001111000000010000000100000000000000011111111100000000000000000000000000101110000000011111000000000001000100000001000000000000000011110000000100010000000000001111",
		"00000000111100000000000000001110001000010000000100000000000000010000000111110001000011110000000000001110000000000000111100000000000000000001111000000000000011110000000000010000000000000001000000000001000000000000000000000000000100000000000000010000000000001111111111100000000000010000000011111111111000000000000111100000000100000000000000000000000000001111000000000000000000011111000000000000111000000000111100000000000000011110000000011110000000010000000000000000000000000000000011110000000100010000000100010000",
		"00000000000000000000000000000000000100000000000100000000111100010000000000000010000011110000000000001111000000010000000000000000000000000000111000000000000000000000000100000000000000000000000000000001000000000000000000000000000100000000000000000000000000001111111111100000000100000000000011111111111100000001000010100000000100000000000000000000000000001111000100000000000000010000000000011111111100000001111100000000000000011110000000001111000000000000000100000000000000010000000000000001000100001111000000010000",
		"00000000000000001111000000000001000011100000000000010000000000000000000011110000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001111000000000001000000000000000000000000000100000000000100000001000000000000000000000000000000000001000000001111000000000000000011000000000000000000000000000000000000000000000100010000000000000000000000011111000011110000000000011111000000001110000000001111000000000001000100000001000000010000000011110000000100000000000000000000",
		"00000000000000000000000000000000000011010001000000010000000000010000000011110000000000000000000000000000111100000000000000000000000111110001000000000000000100000000000100000000000000000000000000000001000000000000000000001111000000000000000000000000000000001110000000000000000000000000000011110000000000000000000011010000000000000000000000010000000000000000000100000000000000000000111100001111000000000000000000100000000000001111000100000000000100000001000000000000000000010000000000000000000000000000000111110000",
		"00000001000000000000000000000000000011110000000100010000000000010000000100000000000000010000000000000000000000000001000000000001000100000000000000000000001011110001000100000000000000000000000000000001000000000000000000010000000000000000000000000000000000001111000000000001000100000001000011110000111100000000000000000000000100000000000000000000000000001111000100000000000000010000111111110000000000000001111100010000000000001110000100000000000000000000000100000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000100000000000000010000000000000000000000000000000000010010000000000000000000000000000000000000000100000000000000000000001011110000000100010001000100000000000000000000000000000000000000000000000000000000111100001110000000000000000000000001000000010000111111110000111100001111000000000000000000000000000011110000000000001111000011110000000000100000111000000000000000000001000000000000000000000000000100000000000000000000000000000000000000010000000000001111000000000000000000000000",
		"00000000111100000000000000000000000100000000000000010000111100000000000000000000000000000000111100000000000000010000000000000000000000001111000000000000000100000000000000010000000000010000000000000000111100000000000100000000000000000001000000001111000100000000000000000010000000010000111100001110000000001110000000000000000000000000000000000000000000000000000011100000000000110000000011100000000100000001000000010000000000000001000000001111111100010001000100011111000000000001000000011111000000000000000000000000",
		"00000000000000000000000000000000001000000000000100010000111100000001000100010000000111110000111000000000000000000000000000000001000000000000111100000000001000000000000100000001000100000000000000000001111000000000000000000001000000000001000000000000000011110000000011110010000100010000000000001110000000001110000000001111000000000000000011110000000000000000000000000000000000000001000011110000000000000000000000000000000000000000000000000000000000000001000100000000000000000001000000011111000000000000000000000000",
		"11110000000000000000000000001111000000010000000100100000000000000000000000000000000000000010000000010000000000001111000000000001000000000000111100000000000111110000000100010000000000010000000000000000000000000001000000000001000000000000000000001110000000000001111100000001000100001111000000001101000000001110000000001111000000001111000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000001000000000000000000000001000100000000000000001111000011110001",
		"00000000000000000000000000000000000000010001000000010000000000000000000000000000000000000011000000010000000000000000000000000001000000000000111100000000000000000000000000010000000000010000000000000000111100000001000000000001000100000000000000011111000100000000000000000001000011111110000011110000000000000000111100000000000000001110000000010000000100001111111100000000000000010000000000000000000100000000111100000001000100000000000000000000000000000001000000010000000000010000010000001111000000000000000000000001",
		"00000000000000001111000111111111000000010001000000000001000000000000000000000000000000000010000100000000000000000000000100000001000000000000111100000000000000000001000000000000000000010000000000001111000011110001000000000000000100000000111000011111000000000000000000000000000100000000000011110000000011110000111100001111000000001110111100000000000000011111111011110000000000000000000000000000000100010000000000000000000011110000000000000000000000010001000000000001000000000001000100011111000000010000000000000000",
		"00000000000000000000000100000000000000000001000011110000000000000000000000000000000000000010000100000001000000001111000000000001000000000000111100000000000000000001000000000000000100100000000000000000111111110010111100000000000100000000111100010000000000000000000000000000000000001111000011111111000000000000111100000000000000001111111000010001111100000000111111110000000000010000000000000000000100100000000000000000000000000000000000000000000000000000000000000001000100000000000100001110000000000001000000000000",
		"00011111111100000000000000000000000000000000000000000000000000100000000000000000000000010000001000000000000000000000000000000001000000000010000000000000000000000001000000001111000100010000000011101110000011110010111100001111000100000000000000100000111100010000111100001110000000000000000000000000111100000000000000010000111100001111000000000001000000010001111100000001111100000000000000000000000100100000000100001111000011110000000000100001000000011111000000000000000000000000000000010000000000000000111100000010",
		"00100000111100000001000111110000111111110000000000000000111000010000000000000000000000000011000000000000000011110000000011110010000011110001111100000000000000010000000000000000000100000001000011111111000111100010110100000000000111110001000000011111111100001111111000001110000000000000000000001111000000001101000000000000111100001111000000000010000000010000000000000001000000000000000111110000000100100000000000010000000011100000111100100010001000011110000100000000000000000001000000000000000000000000000000010001",
		"00010000111100000000000000001111111100000000000100000000111100100000000000000000000000000010000100000000111100000000000011110010000011110001000100000000000000100010000000000000000000000000000000001111000111110001111000011111001000000000000000001111111100001110111000001110000000000000000000001111000000011111000000000000111100000000000000000001000000010000000000000000000000000000000000000000000100011111000000010000000011110000000000100001000000001110000000000000000000000001000000000000000000000000111000010001",
		"00010000000000000000000000001111000000000000000000010010000000010000000000000000000000000000000100000000000011110000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000100000001000000000000000100000000000000000000111100011111000000000000000000000000000000001111000000001111000100000000000000000000000000000001000100000000000000001111000000000000000100000000000100100000000000010000111100010000111100010000000000000000000100000000000000000000000000010000000000010000000000000000",
		"00010000000000000000111100000000000000011110000000010001111100010000111111110001000000000000001000000010000100000000000000010000000000000001111100011111000000010000000000011111000000100000111100011110000100000000000000000000000100000000000111111111000000010001001000000001000011110000000000000000000000011110000100000000000000011111111100000000001000001111000100011111000000000000000000000000000100010000000000010000111100010001111100000000000000000000000000010010000000010000000000010000000100000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000100000000000100100000000100010000111111110000000100000000000100000000000000001111000000000000000100010000000000010001000000000000000000010000000011110000000000001111000000000000000000000000000000010001000100000000111100010000000000000000000011100001000000000000000000000001000000001111000000000000000000000010000000000001000000000000000000000000000100010000000000000000000000100000111011110000000000000000000000000000000100000000000100000001000000000000111100001111111111110001000000000000000011111111",
		"11110000111100000000000000001111000100000000000011110000000100000000000100000000000000000000000000001111000011110001000000000000000000000000000000000000000100000000000000000000111100000000000000000000000000010000000000000000000000010000000000000000000011110000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000001111000000000000111100000000111100000000000100000000000111110000000000000000000100000000000000000000111111110001000000000000000000000000",
		"00000000000011110000111100010000000000000000111100000000000000000001000011110000000011111111000111110000001000000000000000010001000000000000000100000000111100000000000000001111111100001111111100010000000100000000000000010000000100000000000000000000000000000000000100000000111100001111000000000000000000001111000000000000000000010000000000001111000000000000000000011111000000011111111100100001000000000000111100000000000000010000000011100000000011110000000100000000000000000000111100000000000000010000111011111111",
		"00001111000000011111000000010000000000000001000000010000000100000001111111110000111111111111000100001111000100011111000000000000000000000000000000000000111100000001000000001111000000001111000000000000000000000000000000110001000000000001000100010000000000000000000100000000000000001111000100001111111100000000111100000001000000010000111100001110000000000000000000010000001000000000000000110000000000010001111111100000000000000000000011100000000000000000001000000000000000000000111100000000000000100001111111110000",
		"00000000000000000000000000000000000000010000000000000000000000010001000000000000111111111110000000001111000000001111111100000000111111110000000000000000111100000001000000000000000000010000000000000000000000010000000000010000000000000000000100000000000000000000000000000000000000001111000000000000000000001111000000000000000000100000111100011111000000010000000000010000001000000000111100100000000000000001111011110000000011110000111111111111000000000000000111110000000000000000000011100000000000000001000011101111",
		"00000000000000000000000000011111000000010000000000000000000000000000000000000001111011101110000000001111000000001111111100000000000000000001000000000000000000001111000000000000000000100000000000010001000000000000000000000000000000000000000000000000000000001111000000001111000000000000111111110000000011111110000000000000000000100000111000000000000000000000000000010010001000001111000000100001000000010001111100000000000000001111111100001111000000000000000011110000000000000001000011110000000000000000000011110000",
		"00010000000000000000111100000000000000010010000000001110000000000000000000000001111100000000000000000000000000001111000000000000000000000000000000000000111100000000000011110000000000010000000000010010000000000000000000000000000000000001000000000000000000001111000000000000111100010000000000001111111100000000000011100000000000001111111000000000000100011111111100000001001000000000000000010001000000011111000000000001000000000000000000011111000000000000000000000000111100000000000011110000000000001111000000000000",
		"00010000000000010000000000000000000000100001000000010000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000111000010000000000000000000000001111000000000010111100000000000000000000000000000000000000000000000000011111000011110000111100010000000000001111111100000000000011100000000000000000111100000000000000011111000000010000000000000000000100000001000000011111000011110000000000001110000000010000000000000001000000000000000011110000000011110000000000000000000000000000",
		"00000000000000000000000000001111000000000000000000010000000000000000000100000001000000000000000000100000000000010000000000000000000011110000000000000000000000000000000000000000000100010000111111110000000000000000000000000000000100000000000000000000000000001111000000000000111100000000000000000000111100000000000011110000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000011101000000001111000000000000000000000000000000000000000111110000000000001111000000000000",
		"00000000000000000000000000000000000011110001000100000000000000010000000000000001000100000000000000100000000000000000000000000000000011110000111100000001000000000000000000000000000000000000000000000000000000000000000000000000000111110001000000010001000000001111111111110000000000011111000000001111000000001111000000000000000000000000000000000000000000001110000000000000000100000000000000000000000000000000000000000000000000011110000000001111000000000000000000000000000100000001000111100000000011110000000000000000",
		"00010000000000000000000000000000000011100001000000000000000000010001000000000001000000000001000000010000000000000000000111110000000000000000000000000001000000000000000100000000000100000000000000000001000000000000000000000000000100000000000000010001000000001111000000001111000000000000000011101111000000001111111100000000000000000000000000000001000000001110000000000000000100000000000000000000000000000001000000000000000000011111000000000000000100010000000100000000000100000001000011100000000000000000000000000000",
		"00000000000000000000000000000000000011010000000000000000000000010000000000000000000000000000000000010000000000000000000100000000000000000000001000000000000000000001000100000000000000000000111100010010000000000000000000001111000100000001000000000001000000001111000000001110000000010000000000000000000000001111000011110000000000000000000000000000000000001110000011110000000100000000000000000000000000000001000000000000000000000000000011111111000000010000000100000000000000000001000011110000000000000000000000000000",
		"11110000000000000000000000000000000011110000000000010000000000000000000011110000000100000000000000000000000000010000000000000000000000000001001000001111000000010000000000000001001000010000000000000001000000000000000000001111000000000000000000000000000000000000000000001111000000010000000011110000000000000000000000000000000000000000000000000000000100001111000111110000000000000000000000000000000000000001000000000000111100000000000000000000000000010000000000000000000000000000000011110000000000000000000000000000",
		"00000000000000010000000000000000000000000000000000010000000000000000000000000000000000001111000000000000000000000000000100000000000000000000000000000000000000000000000000000001001000100000000000000001000000001111000000000000000000000000000100000000000000000000000000000000000100000000000011110000000000000000000000010000000100000000000000000000000100000000001000000001000000000000111100000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000010000000000010000000000000000000000010000000000000000000011110000000000000000000000000000000000000000000000000000000000000000111100000000000100000000000100000000001000100000000000000000111100000000000000000000000000000000111100000000000000001111000000000000000000010000000011110000000000001111000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000001111000000010000000000000000000000000001000000000000000000000000000000000000",
		"00000000000000010001000000000000000100010000000000010000000000000000000000000000000000000000111100000000000000000000000100000000000011110000000000001111000000000000000100000001000100010000000000010000000000000000000000000000000000000000111100000000000000000000000000000000000100010000000000000000000000001111000000000000000000001111000000000000000000000000000011110000000000000000000000000000000000000000000000000000111100000001000000000000000000010000000000010000000000000001000000010000000000000000000000000000",
		"00000000000000000000000000000000001000000000001000000000111100000000000000000001000100000001111100000000000000000000000000000000000011110000111100000000000100000000000100000001001000010000000000000000111100000000000000000001111100010000000000000000000100000000000000000001000100010000000000000000000100000000000100000000000000000000000000001111000000000000000011110000000000000001000011100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000111100010000000000000000",
		"00000000000000000000000000001111001000000000000000000000000000010000000000000001000000000010000000000000000000000000000000000000000011110000111000000000000000000001000000000000000100010000000000000000111100000000000000000010111100000000000000000000000000000000000000000000001000001111000000000000000100000000000000001111000000010000000000000000000000000000000011110000111100010001000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000010000000011110000",
		"11111111000000000000111100001111001000000000000000010000000000000000000000000000000011110001000000000000111100000000000000000001000000000000111000000001000100000000000100000001000100000001000000011111111100000001000000000010000000000000000000001111000000000001000000000000000100001111000011110000000000000000000000100000000000000000000011110001000000000001000000000000111100110000000011100000000000000000000000010000000000000000000000000000000000000000000000000000111100000000001000001111111100010000000000000001",
		"00001111000000000000000000000000001000000000000100001111000000000000000000000000000000000001000000000000000000000000000000000000000000000000111000000001000000000000000000000000000000010000000000001111000100000001000000000000000100000000111000001111000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000001000100000000000100000000000000000000000000000000000000000000000100001111000000000000000011110000",
		"00000000111100000000000000010000000000010000000000000000000000000000000100000000000000000010000000001111000000001111000000000001000000000000111000000001000100000000000000000000000100000001000000001111000000010010000000000000000100001111111000001111000100000000111111110000000000001111000000000000000000000001000000010000000000010000000000000000000000010000111100000000000000010000000000000000000000000010000000000000000000000000000000000000000000011111000100000000000000001111000100001111000000000000000000000000",
		"00000000111100001110111100010001000000001111000000000000000000010000000000000001111100000000000000000000000000000000000000000001111100000000111100000000000000000001111111110000000100000000000000001111000000010010111100000001000100000000000000000000000100000000000000000000000100001111000000000000111100000000000000010001111100010000000000000000000000100000111100010000000000001111000000000000000000000000000000000000000011110001000000000000000000001110000000000000111100011111000100000000000000000000111000010001",
		"00011111111111111111000000000000111111100000000011110000000000010000000000000001000000000010000100000000000011110001000000000010000000000000000000000000000100000001000000000000000000010000000000001111000100000010111100000001000100000000000000011111111100000000000000001111000100000000000000001111000000001101000000010001111100010000000100000001000000100000000000010000111100000000000011110000000100100000000000000000000011110001111100010001000100001101000000000000000000000000000000000000000100000000111100000010",
		"00101111000000000000000000000000000000000000000000000000111100100000000000000001000000000001000000000000000000000000000000000001000111110000000100000000000000000010000000000000000000100001000011111111000011110000111000000000001100000001000000000000111100000000000000001111000000010000000000001111000100001110000000000000111100000000000000000001000100101110000000000000000000000000000100000001000000010000000000010000000000000000000000000000000000011110000100000000000000000000000000010000000100001111111100000001",
		"00101111000100000000111100001110000000001111000000010001111100101111000011110001000000001111000100000001000100000010000000010000000000000010000000001111000000010000000000010000000000010000111000010000000100000000000000001111000100000000000011111111000000010000000100000001000000000000000000000000000011111111000100000000000000011111000000000000000111110000001000011111000000010000000000000000000100100000000000010000111000010001111100010000000000000000000000010001000000010000000000100000000100010000000111110000",
		"00010000000000000000111000000000000000001111000000010010111000100000000011100001000000000000000100000001000100010001000000010000000000000001111100011111000000010000000000000000000000011111111100000000000011110000000000000000001000000000000111101111000000010001000100010001000011110000000000000000000000011111000111110000000000001111111100000000001000001111001000011111000000000000000000000000000100101111000100000000111100010010111100000000000000000000000000010001000000010000000000010000000100001111000111110000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000111100000000000011110000000000000000111100000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111000000000000111100000000000000010000000000010000111100000000000000001111000000000001000000000000111111110000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000111100000001000000000000000000001111000000000000000000000000000000000000000000000000000000001111000000001111",
		"00000000000000000000000000000000111100000000000000000000000000000000111100000000000000010000000000000001000100000000000000000001000000000000000000000000000000010000000000000000000011110000000011110000000000000000000100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000010000111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000001000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000011111111000000000000000000000000111100000000000000000000000000000000000011110001000000000000000100000000000100000000000000100000111000000000000000000000000000011111000000001111000000000000000000010000000000010000000000000000000000010000000000000000000100000010111111110000000000001111000000000000000011110000000000010000000000001110111100000000111100010000000000000000000000010000000000000010000011110000000000000000000111100000000000000000000100000000000000000000111100100001000000001111000000001110",
		"00100000000100000000111100000000000000000000111100000000000000000001000000000000111111110000000011110000000000000000000000000000111000000000000000000000000000000000000000001111111100000000111100000000000000000000000000000000000000000000000000000000000011110000000100000000111100000000000111110000000000001111000111100000000000000000111100001111000000000000111100010000000100000000111100100001000100010000111100000001000000000000000011110000000000000000000000000000000000000000111100100000000000010000111111111111",
		"00010000000000001111000000010000111100010000000100000000000000000010000000000000111111110001000000001110000000011110000000000000111100010000001000000000000000000001000000000000000100010000000000000000111100010000111000100000000000000000000000011111000000001111000111100000000000001111000000000000000000000000000000001111000000000000111100001111000100011111111100000000001000001111111100100000000100100001000000000001000011110000111100001111000000000000000011111111000000000000111100010000111100010001111111110000",
		"00000000000000001111111100001111000000101111000000000000000100100001000000000000110111111111000000001110000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000010000000000000001000000000000000000001110000011110000000000000000000000010000000000000000000000010000000000010000111100000000000000011111000000000001001000000000111100010000000000000001111100000010000000000000000011111111000000000000000011110000000000000000000000000000111100000000111100001111",
		"00000000000000000000111100000000000000010000000000001111000100100000000000010000111011111101000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000001111000000000000000000000000111100000000000011110000000000000000000000001111111100000000000000000000111100000010001000000000111100010000000000010000000000000001000000001111111100011111000000010000000011110000111100000001000000000000000000000000000000000000",
		"00000000000000000000000000000001000000100000000100000000000000000000000000010000111100000000000000000000000011110000000000000000000000000000000000000000111100000000000000000000000100010000000000000000000000000000000000010000111100000001000000010000000000001111000000000000111100010000111100000000000000000000000000000000000000001111111111110000000000010000111100000001000100000000000000000001000100000000000000000001000000001110000000001110000000010001000100000000000000000000000000000000111111110000000000000000",
		"00000000000000000000000000010000000000010001000000000000000000000001000000100001000000010000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000001111000000000000000000000000000000000000000000000001000000010000000000001110111100000000111100010000111100000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000001000000010000000000000010000100011110000000011110000000100000000000000000000000000001000000000000111111111111000000010000",
		"00000000000000000000000000010000000000000000000000000000000000000000000000010000000000001111000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000010000000000001110000011110000111100010000000000000000111100000000111100010001000000000000000000000000000000001111111100000000000000000000000000000001111100000001111100000000000000011111000000000000000000011111000100000000000000000000000011100000000000000000000000000000",
		"00010001000111110000000000000001000011100000000100000000000000000000000000000000000000000000000000010000000100001111000000000000000000000000000000000001000000000000000011110000111100000001000011110000000000000000000100000000000000000000111100000001000000000000000000001111000000010000000000000000000000000000111100000000000000000000000000000001000000001110000000000000000000000001000100000000111100000001000000000000000000011111000000000000000000010000000000001111000000000000000011100000000000000000000000000000",
		"00000000000100000000000000000000000011010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000010001000000000000000000000000000000000000000000000000111100000001111100001111000000001110000000100000000011111111000000000000000000000000000000000000000000000000000000001110000011110000000000000001000100000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000011110000000011110000000000000000",
		"11110001000000000000000000000000000011010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000001000100000001000000000001000000000000000000000000000000001111000000000000000000000001000000000000000000001110000000010000000000001111000000000000000000100000000100000001111100000000000000001111000000000000000000000000000000000000000000000000000000000001000000000000000011110000000100011111000000000000000000000000000011110000000000000000000000000000",
		"11100001000000000001000011110000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000001000000000000000000001111000000010000000000000001000000000000000000001110000000010001000000000000000100000000000000010000000100000001000000000000000000000000000100000000000000000000000000000000111100000000000000000000000000000000000000000000000100001111000100000000000000000000000011110000000000000000000000000000",
		"11110001000000000000000000000000000000000000000000010000000000010000000000000000000000001111000000000000000000000001000100000000000011110000000000000000000000010000000100000000000100000000000000010001000000000000000000001111000000000000000000000001000000000000000000000000000000100000000000000000000100000000000000010000000000000000000000000000000011110000000100000000000000000000000000000001000000000000000000010010000000000001000011110000000000000000000000010001000000000001000011110000000000000000000000000001",
		"00000001000000010000000000000000000100010000000000000000000000000000000000000001000000001111000000000000000000000000000100000000000111110000111000000000000000000000000100000000000100010000000000000001000000000000000100001111000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011100000000000001111000000000001000000000001111100000000111100000000000000000000",
		"00000001000000000001000000000000000100000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000111000000000000000000000000000000000000100000000111100000000000000000000000000000000000000000000000000000001000000010000000000000001000000010000000011110000000100000000000000000000000000000001000000000000000000000000000000000000000011110000000011110000000000000000000000000001000000000000000000000000000000001111000000000000000000000000000000000001000011110000000000000001",
		"11110000000000010001000000000000000100000001000000000000000000010000000000010000000000000000000000000000000000000000000000000000000111110000110100000001000000000000000000000000000000000000000000000001000000000000000000000000000000000001000100000001000000010000000000000001000000010000000000000001000100000000000000000000000000000001000000000000000000000001000000000000000000000000000011101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000010",
		"00000000000000010001000000001111000000000000000000010000000000010000000000010000000000000000000000000000000000000000000000000000000011110000111000000000000000000000111100000000001000000000000000000000111000000000000000000001000000000000000000000001000000001111000000000000000000011111000000001111000100001111000011110000000000000001000100000000000000000001000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000011111111100000001000000000000",
		"00000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000100000000000000010000000000000000000000000000111000000001000000000000000000000001001000000000111100000000111000000000000000000001000000001111000000000001000000000000000011110000000100010000000000000000000000001111000011110000000000000010000100000000000000000001000011110000000000000000000011100000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001",
		"11110000000000000000000000000000000000000000000000000000000000000000000000010000111100000000000000000000000000010000000000010000000000001111111100000000000000010000000000000001001000000000000000000000000000000001000000000001000000000000000000000000000000000001000000000001000100010000111100011111000000000000000000000000000000010001000011110000000000000000000011110000000000000000000000000000000000000000000000000000000000001111000000000001000000000000000000000000000000000000000000011111111100000000000000000001",
		"11110000111100000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000001111000000000000111100010000000000000000000000010000000000000000001000000000000000000000000000000001000000000000000100001111000000000000000100000000000000000000001000000000111100000000000000000001000011110001000000000000000000000000000100000000111000000000000000000000000000000000000100000001000000000000000011110000111100000000111100001110000000000000000000000000000100011111000011110000000000000000",
		"00000000111100010000000000000000000000000000000000000000000000000000000000010000111000000000000000000000000011110000000100001111000000000001000000000001000100000000000000000001001000000001000000000000000011110001000000000000000000000000000000001111000000001111000000001111000111111111000000001101000000001110000011100000000000010000000100010000000100010000111000000000000000010000000011111111000100000001000000011111111111110000111100000000000000001111000000000000000000010000001100000000000000010000000000000001",
		"00010000000000010000000000000000000000000000000000000000000000000000000000000001111100010000000000000000000011110010000011100001111100000010000000000010000000000000000100000000000000000001000000001111000000000001111100000000000100000000000000011111000000001111000000001111000111110000000000001110000000001110000100000010000000100000000011110000000000000000111000010000111100001111000000001110000100010000000000011110000011110001000000010000000000000000000000000000000000010000001000000000000000010000111100000010",
		"00101110000000100000111100001111000000001111000000000000111100011110000000000000000100010000000000100000000011110010000011110001000000000000000000000000000100000001000000000001000000010010000100001110001000000001111100000000001000000001000000011111000011110000000000000000000000000000000000000000000100001110000000000000111000100000001000000000000000000000000000000000000000010000000000000000000000010000001000010000111111110000000000000000000100011110000000000000111100000000000000001111000100010000000111110010",
		"00010000000000010000111100000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000011110000000000000000000100000000000000000000000011110000000100000000000000001111000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000011110000000000000000000100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000001111000000000000111100000000000011110000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000100010000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100010000000000000000111100000000000000000000000000000000000000000000000000000000000000010000000100000000000100000000",
		"00010000000000000000000000010000000000000000000000000000000000000000000000011111111100000001000100000000000000010000000000000000000000000000000100000000111100000000111111111111000011111111111100000000111100000001000000000000000011110001000000000000111100000000000000010000000000000001000000000000000000000001111100000000111111110000111100000000000100010000000000000000000011110000000000000000000000011111000011110000000100000001000000000000000000000001111100000000000000000000000000000000111100000001000000000001",
		"00010000000100001111000000001111000011100000000000010001000000010001000000011111000000000010111100000000000000000000000100000000000000010000111100000000000000000000000011111111111111111111111111110001111100000001000000000001111000010010111000000001111000001111000011110000111100000000111100000001000000000000000000000000000000010000000011110000000000001110111000010000000000000001111100010000000000000000111100010000000000001110000011110000000000000001000100000000111100000000111100000001111000011111111100001111",
		"00000000000000000000000000000000000000000000000000010000000000000000000000010000000100000000000000000000000100000000000000000000000000000001000000000000000000010000000000000000000000001111000000000000000000000000000100000000000000000000111100000001000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000111100000000000100000000000000000001000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00100000000000000000000000010000000000000000111100000000000000000001000000010000000000000001000011110000001000000000000000001111000000100000111100000000000000000000000100000000000000001111000000000000000000010000111100010000000000000001000000000000000011110000000100000001111100000000000000000000000100000000000011110000000000000000000000011111111100010000000000000001000100000000000000010001000000000000000000000001000000000000000011110000000000000000000000000000000000000001000000100000000000010000000000001111",
		"00000000000100000000111100000000000000000000111100001111000000000010000000000000111111110000000011100000000000000001000000000000111100000000000000000000000011110000000000000000000000000000000000001111000000010000111100000000000000000000111100010000000011110000001011010001111100000000000000000001000000000000000011110000000000010000111100000000000000000000000011110000000100000000111000000000000000010001111100000001000000000000000011110000000000000000000000000000000000000000111100010001000000010000000000001110",
		"00010000000000000000111100000000000000010000000100001111000000000001000000100000111000000000000000001111000100100000000000000000000000010000000100000000000100000001000000000000001000100000111100000000000000010000111000000000000000000000000000000000000100000000000111100000000000001111000000000000000000000000000111100000000000011111111100001111000100010000000000000000001000010000111000000000000000000010000000000001000000000000000000000000000000010000000011110000000011110000111100000000000000000000111100000000",
		"00000000000000000000111100000000000000000000000000001111000000010000000000010001111111111111000000000000000000010000111100000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000111100000000000000000010111100010001000100001111000011110000000000000000000000000000001000000001000000000000000000000000111100000000000000001111111100000001001000000000000000000000000000000001000000000001000000001111000000001111000100010000000000000000111100000001111100010000111100000000000000001111",
		"00000000000000000000000000000000000000010000000000001111000100010000000000000000111000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000111100000001000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000001111111100000000000100011111111100000001001000000000000000000000000000010001000000000000000000000000000000001111000000100000000011110000000000000000000000010000000000010000000000000000",
		"00000000000011110000000000000000000000010000000000001111000000010000000000000000111100000000000000000001000011110001000000000000000000000000000000000000000000000000000000000001000000010000000000000000000100000000000000000000000000000001000000000000000000000000111100000000111100011111000000000000000000000000000000000000000000001111000000000000000000001111000000000000000100000000000000000000000000000000000000000000000000001110000000011110000000010000000000001111000000000001000000000000000000001111111100000000",
		"00010000000000000000000000000000111100000000000000010000000000000000111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111100010000000000001110000000000000111100000000000000000000000000000000000000000000000000001111000000000000000000001110000000000000000000000000000000000000000000010000000011110000000000000000000000001111000000010000000000000000000000000000000000000000000000001111000000000000",
		"00010000000000000000000000000000000000000000000100000000000000001111000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000001111000000000000000000010000111100000000111000000000000000001111000011110000000000000000000000000000000000000000000000010001000011110000000000000000000000001110111100001111000000000000000000000000111100000001000011110000000000000000111100000000000000010000000000000000000000000000000000000000000000000000000000000001",
		"00000001000000000000000000000000000011100000000100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000010001111111110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001110000000000000000000000000000000000000111100000000000000000001000000000000111100000000000000000000000000000000000000001111000011110000000000000000000000000000",
		"00000000000100000000000000000001000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000111100000000000000000000000100000000000000000000000000000001000000000000000000000000000000010001000000000000000000000000000000010000000000000001111100000000000000000000000011110000000000000000000000000000111100000000000000000001000000000000111111110000000000000000000000000000000000000000000011110000000000000000000011110000",
		"11100000000000000001000000000000000011110000111100001111000000000001000000010000000000000000111100000001000000001111000000000000000000000000000100000000000000000000000000000000000011110000111100010000000000000000000100000000000000000001000000000001000000000000000000001111000000010000000000000000000000000000000000100000000000000001000000000000111100000000000011110000000011110000000000000000111111110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000",
		"11100000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000011111000000010000000000000000000000000000000000001111000000010001000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000000000000000000000000000000000000000000010000000011110000000000000000000011110001",
		"11110001000000000000000000000000000100010000000000000000000000010000000000000000000000011111000011110001111100000000000000000000000000000000111100000000000100000000000000010000000000000000000000010000000000000001000000001111000000000000000000000001000000000000000000000000000000100000111100000000000100000000111100000000000000000001000000000000000000000001000100000000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000001000010000000011110000111100000000000000000001",
		"00000000000000010000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000011110000000000000000000011110000111100000000000100000000111100001111000000000000000000000000000000000000000000001111000000000000000100000001000000000000000000000000000000110000000000010000000100000000000011110001000000000001000000000000000100000000000000000000000000000000000100000000000000000000000000000001000011110000000000000000000000011111000000000000000100000000111111110000111100000000000000000001",
		"00000001000000100000000000000000000000010000000000000000000100000000000000000000000100010000000000000000000000000000000100000000000000000000111100000000000000000000000000000000000111110000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000010000001000000001000011110001000100000000000000000000000100000001000000001111000000000001000011110000000000000000000000000000000011110000000000000000000000000000000000000001000100000000000000000000000000000000000000000001",
		"00000000000000000001000000001111000000000000000000000000000100000000000000000000000000000001000000000000000000000000000100000000000011110000111100000000000000000000111100000000001000000000111100000001000000000000000000000001000000000000000000000000000100010000000011110000000000000000000000010000001000000000000011110000000000000000000000000000000100000001000000000000000000000000000111100000000000000001000100000000000011111111000000000000000000000000000100000000000000000000000000000000000000000000000000000001",
		"00000001000000010001000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000001100000000000000000001111100000001000000000001000000010000000000010000000000000000000000000000000100001111000000011111000100001111000011110001000000000000000000000000000100000001000000000000000000000000000111000000000000000000000100000000000100000000000000000000000000000000000000000000000100000000000000011111000000000000000000000010",
		"00000000000000000000000000000000000000000000000100000000000000000001000000000000111100000000000100000000000000000000000000000000000000000000000000000001000000000000111100010000001000000000111100000000111100000000111100000010000000000000000000000001000000000000000000000001001000000000000000011110000100000000000011100000000000010010000000000000000000000000000111110000000000000000000011100000000000000000000100000000000000001111000000000001000011111111000000000000000000000000000100001111000000000000000000000010",
		"00000000000100000001000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000001111000000000000000000010000111100000001001000000001000000000000000000000000111100000000000000000000000000000000000000000000000000000000000100000000111100010000000100000000000011110000000000000000000100000000000000000000000000000000000000000000000111110000000000000000001000000000000000001111000000000010000000000000000000000000000000000000000100001110000000000000000000000010",
		"00000000000000000000000000000000000000000000000000000000000111110000000000010000000000000000000000000000000000000000000000000000111100010000000100000000000000010000000000000000001111110000000000000000000000000000111100000000000000000000000000000000000000000000000100001111001100000000111100001111000000000000000011010001000000010000000100000000000000000000111100000001000000000000000011110000000000000000000000000000000011110000000000010001111100001110000000001111000000000000000000011111000000000000000000000000",
		"00000000111100000000000011110000000011110000000011110000000000000001000000100000000000010000000000000000111100000000000000001110000000000000000000000000000000010000000000000001001000000001000000000000000000000010000011110000000100000000000000010000000011110000000000001110001011110000000000001111000000001111000011100001000000000000000000000000000100000001111100000001000000000000000100001111000000000001000000001110111111100000000000000001000000001110000000000000000100010000000000000000000000010001111111110000",
		"00000001000000000001000000000000111111111111000000000000000000000000111100010000000000011111000000010001111100000000000000000000000000000001000000000000000000010000000000000010000000000000000000000000000000000000000011110000000111110000000000101111111111110000000000001111000011100000000100001111000000000000000000000000000000001111000000000000000000000000111000000001000000000000000000000000001000000000000000001110111111110000000000001111000000001110111100000001000000000000000100010000000000010000000000000000",
		"00011111111100000001000011100000000000001111001000000000111000011111000000000000001000000000111100010001111100000000000000000000000000000000111100000000000100010001000100000011000000000000000100000000000111100000111000001110000100000001000000010000000000001111000000001111111100000000000000010000000000000000000000001111111100000000000100000000000011110000111100000000000000000000000000000000000100001111000000001111000011111111111100000000000000001110000000000000111100000000000100000000000000000000001000000000",
		"00010000000000000000000000000000000000000000000100000001000000000000000000000000000000000001000000000000000000000000000011110001000000010000000000000000000000000000000011100000000100000000000111111111000000010001111100010000000100000000000000001111111100000000111100000000000100000000000011111101000000001111000100000000111100000000000100000010000000010000000000000001000000000000000111101111000000010000000100000000000000000001000000100010000000000000000100000000000000000001000100000000000000000000000000000000",
		"00000000000000000000111100000000000000001111000000000000000000000000000000000000000000000000000000000000000111110000111100000000000000000000000000000000000000000000000011110001000100000000000000000000000100010000000000000000000000000000000000000000000100010000000000000000000000000000000100000000000000000000000100000000000000000000000000000000111100000000000100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00010000111011110000111000001111000000100000000100100001111000000000000100001110000000001111000000011111001000010000000000001110111100000001001011111110000100000010000000000001000100001111000011101111000111110000000000000000000000010000000000000000000100011110001011100001000000001111111000100001001011100010000011110000000000000000111000100000000111110000111000010000000100000010111100001111000100000000111100000000000000000000000011111111111100100010000100000001000111110000000100000000001000010001000011111111",
		"00001111001000000000000000001111000011110000000000001111000000000000000000000000000100000010111100000000000100000000000000000000000000000000111000000000000000010000000011110000000011110000111111100001000000000000000000000000111100000001111100000001000000010000000111110000000000000000000000011111000000000000000011100000000000000000000011110000111100001111000000010000000000000001111100000000000000000001000000000000000100001110000000000000000000000000000000010000111111111111111100000000000000010000000000100000",
		"00000000000000000000000000000000000000000000000100000000000000000000111100000000000000000001000000000000000111110000000000010000000000000000000100000000000000000000000000000000000000010000000011110000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000011100000000000000000000000010000000000000000000000000000000100000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000001000000000000",
		"00010001000000000000000000001111000000000001000000000000000000000001000000010000111100000001000011110000000100001111000000000000000100010000111100000001000000000000000000000000000000001111000000000000000000010000000000000000000000000000000000000000000000000000001011110000111100000000000000000000000100000000000011110001000100000000000000000000000000000000000011110000000011110001000000010000000100000000000011110001000000001111000000000000000100010000000000010000000000000000000000100010000000000000000011111111",
		"00000000000000000000000000000000000000000000000000001111000000000010000000000000111000000000000011110000000000000000000100000001000000000000000000000000000100000001000000000000000000001111111000000000000000101111000000000000000000010000000000011111000011110000001011110000111111100000000000000000000000000000000000000000000100011111000000000000000100000000000000000000000100000000111100000000000000000000111100000000000000000000000000000000000100000000000000000001111100000000111000000001000000010000111111101111",
		"00000000000000000000000000000000111100000000000000000000000011110001000000000001111000000000000000000000000000010000000000000000000000000000000000000000000100000010000000000000000000010000111100000000000000000000111100000000111100000001000000000000000000000000000000000000111100000000000000001111000100000000000011100000000000011111000000011111000000000000000011110000001000010000000000000000000000000001000000000000000111110000000000000000000000100000000000000000000011110000111000000000111100000000111100001111",
		"00000000000000000000000011110000000000000000000000000000000000000001000000010000111100000000000000000000000000010000000100000000000000000000000000000000000000000000000100000000000100010000000000000000000000000000000000000000111100000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000111100000000000011110000000000010000111100000000000000000001000000010000111100000000000000001111",
		"00000000000000000000000000000000000000000000000000010000000000000000000000000000111000000000000011110001000000000000000000000000000000000000000000000000000100000000000000000000000000000000111100000000000000000000000000000000111100000001000000000000000000001111111100000000000011110000000000000000000000010000000000000000000000000000000000000000000100000000111100000000001000000000000000000000000000010001000000000000000011110000111100001111000000010000000000010000000000000000000000010000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000111100001111000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000010000000000000001000000000000000000000000000000001111111100000000111100000000000000000001000100000000000000000000000000000000000011111111000011110000000011110000000011110000000000000000000000000000000000001111000000011111000000100000000000000000000000000001000000010000000011111111000000000000",
		"00010000000000000000000000000000000000010000000000011111000000001111000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000111100011111000000000000000000000000000000000000000000000000000000000000000000000001000111110000000000000000000000001110000000001111000011110000000000000000000000010000000000000000000000001111000000011111000000010000000000000000000000000000000000000000000000001111000000001111",
		"00000000000000000000000000010000000000000000000100000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000111000000000000000000000000000001111111100000000111111110000000000000000000000000000000000000000111111110000000000000000111111110000000000000000000000000000000100000000000000010010000100000000000000000000000000001110000000000000000000000000000000000000111100000000111100000001000000001111000000000000000000000000111100000000000011111111000000000000000000001111000000000000",
		"00000000000000000000000100000000000011100000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000111111110000000000000000000000000000000100000000000011110000000000000000000000000000000000000000000000000000000100000000000000010001000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000010000100000000000011100000000000000000000000000000000000001111000000000000000100000000000000000000",
		"00000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000100001111100000000000000000000000000010000000100000000000000000000000000000000000011110000111100001111000011110000000000000001000000010000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000001111100000000000000000001000000000001111111100000000000000000000000000000000100001111000000000000000100000000000011110000",
		"11110000000000000000000000000000000011110000111100000000000000000001000000000000000011110000000000010001111100000000000000000000000000000000000100000000000000000001000000000000111100000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100001111000000001111000000000000000000000000000000000000000011110000000000000000111100000001111100000000000000010010000000000001000000000000000000000000000000000000000000010000000000000000000000000000000011110000",
		"11110000000000000000000000000000000000000000000000000000000000000001000000000000000000001111000000000001000000000000000000000000000000000000000000000000000000000001000000010000111100000000000000010000000000000000000000011110000000010000000000000001000000000000000000001110000000010000000000010000000100000000000000000000000000000001000000001111000000000000000000000000000100000000000000010001000000000000000000000010000000000001000000000000000000000000000000000000000100010000111100000001000000000000000000000000",
		"00000000000000010000000000010000000000010000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001000000000000000000011110000000010000000000000001000000001111000000000000000000010000111100100000000000000001000000000000000000000000000000001111000100000000000000000000000011110000000100010000000000000000000000000000000011110000000100001111000000000000000100000000001000000000111100000001111100000000000000000000",
		"00000001111100000000000000010000000000010000000000000001000000000001000000000000000000010000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000100000000000000000001000000000000000000001111111100010000000000000001000000000000000000000001000000010000111100010000001000000001000011110000000000000001000000000000000100000001000100001111000000000000000011110000000000000000000000000000000000001111000100000000000000000000000100000000000100000000111111110010111100000001000000000000",
		"00000000000000000000000000000000000000010000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000000001000100001111000011110001000000000000000000010000000100000001000011110010000000000000000000000000000100000000000000001111000000000001000111110000000000000001000100000000000000001111000000000000000000001111000000010000000000000000111100000001000000000000000000000000",
		"00000000000000000001000000001111000000000000111100001111000000000000000000011111000000000000000000000000000000001111000100000000000100000000000000000000000000000000000000000000000111110000000000000010000000000001000000000001000000000000111100010000000000000000111111110001000000000000000000000000000100000000000000000000000000000001000000000000000100000001000000000000000000000000000011010000000000000000000100000000000000001111000000000000000100011111000000000000000100000000111100000000000000000000000000010000",
		"00000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000001111000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000100001111000000000001000000000000000000000000000100000000000000000000000000000000000111100000111100000000000100000000000000000000000000000000000100000000000000000000000000000000000000001110000000000000000000000000",
		"00000000000000000000000000001111000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000111100010000000100000000000000000001000000000001000000000001000000000000111100000000000000000000000011110001001000000000000000010000000100001111000011110000000000010000000000000000000000000000000000000000000000000000000111110000000000000001001000000000000000000000000000000000000000000000000000000000000000000000001000001101000000000000000000000000",
		"00000000000000000000000000001111000000000000000000000001000100000000000000000000000000000000000000000000111100000000000000000000000000000000001000000000000000000000111100000000000111110001000000000001000000000000000000000000000000000000000000000000000011110000000000000000001000000000000000000000000100000000000011110000000000000000000000000000000000000000000000000000000000000000000100001111000000000000000100010000111100000000000000000001000000000000000000000001000000000000000000001101000000000000000011110000",
		"00000000000000000000000000000000000011110000000000000000000100000000000000010000111100000000000000000000111100001111000000000000000000010000000000000000000000000001000000000000000100000001000000000000111100000001000000000000000000000000000000000000000011110000000000001110000100000000111100000000000000010000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000100000000000011110000000000000000000000000000000000000000000000010000000000001110000000000000000000000000",
		"00000000000011110000000000000000000011111111000000001111000100000000000100010000000000000000000000000000111000000000000000001110000000010000000100000000000000010001000000000001000111110000000000000000000000000001000000000000000000010000000000001111111100000000000011111111000000000000000000001111000011110000000011100000000000000000000100001111000000000001111100000000000000010001000000000000000011110001000000000000000111100000000000000000111100001111000100001111111100000000000000001111000000010001000011111111",
		"00000000111100000000000111010000111111110000000100000001000000000001000000100000000000000000111100000000111100010000000000001111111100000000000000000000000000100000000000000010000111110000000100000000000011100001111111111101000000000000000000011111111011110000111100001110000000000000000100000000000011100000000011111111000011110000000100000000000000000000111011110001111100000000000000000000000100000000000100011110111100000000000000000000111000001110000000000000000011110000000100001111111100000001000000001111",
		"00000000000000000000000011010000000000000000001100000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000011110010001000000000000111110000000000000001000000001111000100001111000000000000111111110000111100001110000100001111000000001101000000001111000111110000000011100000000100000000000000000000111111100001111100001110000000001110000100000000000100000000000011100000000000010000111100001111000000000000000000000010001011111111000000000000000000000000",
		"00000000000000000000000000000000000100001111000100000000000100000000000000000000000100000001000000000000000011110000000000000001000000000000111100000000000000000000000011110001000100000000000000001111000100010001000000010000000011110000111100001111111100000000000011110000000100000000000011111111000000001111000111110000000000000000000100000010111100000001000100000001000000000000000011110000111100010001000000010000000000000000111100100001000000011111000000000000000000000000000011100001000000010000000000000000",
		"00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000100000000000000000001000111110000000011110000000000010000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000011110000111100000001111100010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
		"00000001000100000000000000000000000011110000000000000000000000000001111100011111111100000001111100000000000100001111000000000000000000010000000100000000000000010000000011110000000011110000111011110001000011110001000100000000000000000001111100000001111100010000000011110000111100000000000000000000000000000000000011100001000011111111111100000000000000000000111100000000000011100000000000000000000100000000000000000000000011111111000000001111000100010000000000000000000011110000111100000000111100010000000000000000",
		"00000000000011110000000000001111000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000100000000000000000000000011111111000000000000000000001111000000000000000000000000000100000000000000000000000000000000",
		"00000000000000000000000100000000111100000010000011111111111100000000000000001111000100000000000011110001000000000000000011110000000100000000111100000000000000000000000111110000000011111111000000000000000000010001000000000000000000000000111100010001000000000000000011110000111100000000111100000000000100000000111100000000000100000000000000000000000011110000000000001111000011110001000000010000000000000000111000000001000100000000000000001110000100010000000100011111111100001111000000100001000000110000000000001111",
		"00000000000000001110000000000000111100000000000000001111000000000010000000000000111000000000000000000000000000000000000100000000000000000000000000000000000000000001000100000000000000011111111000001111000000000000000100000000111000010000000000000000000100000000000100000000111111110001000011110000000000010000000000000000000100100000000000000000000000000000000000000000000100000000000000010001000000010001000000000000000011110000000000000000000000000010000000000000111100000000111100000000111100010000111011100000",
		"00000000000100000000000000000000111100000000000000000000000000000001000100010000111000000000000000000000000000000000000000000000000000001111000100000000000000000000000100000000111100001111111100001111000100001111111100000000111100000001000000000000000000001110000000000000111100000000000000000000000000000000000000000000000000010001111100010000000000001111000000000000001000000001000000000001000000000000000000000000000111110000000111111111000100100000000000000000000011110000111100000000000000001111111000000000",
		"00000000000100000000000000001111000000000000000000000000000000000001000000010000111100000000111100000001111100000000000000000000000100000000000000000001000000000000000011110000000000000000111100000000111100000000000000000000111111110010000000000000000000011111000000001111000011110001111100000000000000000000000000000000000000000001000000000000000000000000000000000000001100000000000000000000000000000000000000001111000000000001000000000000000000010000111100000000000000000000111100000000000000000001000000001111",
		"00000000000100000000000000000000000000011111000100000000000000000000000000001111111111110000000000000000000000000000000000000000000000000001000000000000000000000000000011110000000000000000111100001111000011110000000000000000000000000001111100000000000000001111000000000000000011110000111100000000000000000000000000000000000000000000000000000000000000001111000000001111001000000001000000000000000000000000000000000000000000000001000000001111000000010000111100001111000000000000000000000000000000010001111100001111",
		"00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000011111111000000000000111100000000111100000000000000000000000000000000111100000001000000000000000000000000111100000000000000000000111100000000000000010000000000000000000000000000000000000000000000001110000000001111000000000000000011110000000000000000000000000000000000000000000000011110000000010000000000001111000000000001000000001111000000000000000000000000",
		"00000000000000000000000100000000000000000000000100001111000100000000000000000000000000000000000000000001111000000000000000000000000100000000000000000000000000000000000000000000111100000001000000000000000000000000000000000001000011110000111100000000000000000000000000000000000111110000111100000000000000000000000000010010000000000000000000000000000000001111000000000000000000000000000000000000111100000000000000000001000000011111000000010000000000000000111111110000000000000001000000000000000000000000000000000000",
		"00000000000000000000000100000000000000000000000100000000000000001111000000000000000000000000000000000000111000000000000000000000000100010000111000000000000000000000000000000000000000000001000011110000000011110000000000000000000000000000000000000000000000000000000000000000000100000000000000010001000100000000000000000001000000000000000000000000000000001111000000000000000000000000000011110000000000000000000000000001000000001111000000000000000000000000111100000000000000000000000000010000000000001111000000000000",
		"00000000000000000000000100000000000011110000000100000000000000000000000000000000000000000000000000100000111000000000000000000000000000000000000000000001000000000000000000000000000011110000000011110000000011100000000000000001000100000000000000000000111100000000000000000000000011110000000000000000000111110000111100000000000000000000000000000000111100000000000000000000000000000000000000000001000000010000000000000001000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000",
		"00000000000000000000001000000000000011100000111100000000000000000000000000010000000000000000000000100001111100000000000000000000000000010000000100000000000000000001000000000001000000000000000000000000000000000000000000000001000100000001000000000000111100000000000000000000000011110000000000000000000111110000000000000000000000000000000011110000000000010000111111110001000000000000111100000010000000010000000000000001000100000000000011110000000000000000111100000000000000010000000000010001000011110000000000000000",
		"00000000000000000000000011110000000000000000111000000000000000000001000000010000000000000000000000000001111100010000000000000000000000000000000100000000000000000010000000000000000000000000000000011111000011110001000011110000000000010000000100000000000000000000000000001111000011110000000000100000000100001111000000001111000000000001000000001111000000000000000011100000000000000000111100000001000011110000000000000000000000000000000011110001000100000000111100000000000000010000000000000001000011110000000100000000",
		"00000000000100000000000011110000111100000000111100000000000000000001000000000000111100000000000011110001000000000001000000000000000100010000000000000000000000000001000000000000111111110000000000010000000011110001000000001110111100010000000000000001000000000000000000001101000011110001000000100000000100000000000000001111000000000001000000001110000000010000000000000000000000000000111100010001000011110000000000000000000000000001000011110000000000010000111100000000000000000000000000000001000000000000000000000000",
		"00000000000100000000000000010000000000100000000000000000000100000001000000000000000000000000000011110000000000000000000000000000000100000000000000000000000000000000111100000000000100000000000000010001000000000000000000001101111100000000000000000001000000000000000000000000000011110000000000100000000000000010000000000000000000000001000011110000000000000000000000000000000000000000000000010000000011110000000000000000000000000000000100000000000000000000000000000000000000000000111000000010111100000000000000001111",
		"00000000000000010000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000100000000000011110000000000000000000000000000000000000000111100000000000100000000000000000000000100000000111100001111000000000000000000000001000000000000111100000010000000000000111100100000000000000001000000000000000000000000000011110000000100000001000000000000000000000000000011110000000000000001000000001111000000000000000100000000000000010000000000000000000100000000111100000010000000000000000000001101",
		"00000001000000000000000000000000000000010000000000000000000100000001000000000000000000000000000000000000000000001111000000000000000100010000000000000001000000001111000000000000000011110000000000000001000000000000111100000001000000000000111000000001000011110000111111110001000000000000111100010000000000000000000000010000000000000000000000001111000011110000000000000000000000000000000011110000000000000001000000000000000000000000000000000000000100000000000000000000000000000000111100000010000000000001000000001101",
		"00000000000011110000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000010000000100100000001000000001000000001111000000000000000000000000000100000000000000000000000000000001111100000000000000000000000100000000000000000000000100000000000000010000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000011100000111100000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000001110",
		"00000001000011110000000000000000111111110000111100000001000100000000000000000000000000000000000000000000000000000000000000010000000100010001001000000000000000001111000000000000000100000000000000000001000000000000000011110001000000000000111100010000000000000000000000000000000100000000111100010001000100000000000000000000000000000000000000000000000011110000000100000000000000000000111111100000000000000000000000000000000000001111000000000000000000000000000000010000000000000000000100001100000000000000000100001101",
		"00000001000011100000000000000000000011110000000000000000000000000000000000001111000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000001111000000000001111100000000000000000001000000000000111100000000000000000000000011110000000000000000000000000000000100000000000011111111000000000000000000001111000000000000000100000000000000000000111100000000000000000000000000000000000000001111000000000000000000000000000000010000000000000001000100001100000000000000000000001101",
		"00000000000011100000000000001111000000000000111100000000000000000000000000000000000000010000000000000000000000011111000000000000000000000000000100000000000000000000000000000000000000000000000000000000111100000001000000000000000000000000000000000000000011110000000000001111000100000000000000000000000000001111000011110000000011110000000100000000000000000000000000000000000000000000000000001111000000000000000000010000111100000000000000010001000000000000000000000001000000000000000000001101000000000000000000001101",
		"00000000000011110000000000001111000011110000111000000000000100000000000000000000111100000000000000000000110100001111000000000000000000010001000000000000000000000000000000000000000011110000000000000001000000000010000000010000111100000000000000000000000011110000111100001111000000000000000000000000000000010000000011110000000000000000000011110000000000000000000000000001000000000000000000000000111100000000000000000000000011111111000000000000000000000000000000000000000000010000000000001111000000010000000000001110",
		"00000000000111110000000000001111000111110000111100000000000000000000000100000000000000010000111111110000000000001111000000011111000000000000000000000001000100000000000100000000000011110001000000000000000011110000000000000000000000000000000000010000000000000000111100001110000000000000000000000000000000001111000011100000000000000000000100000000000000000000000000000000000000000001111100000000000011110001000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000010000000000001101",
		"00010000000011110000000011100000000011111111000000010001000100000000000100011111000100010000000000000000000000000000111100000000000000000000000100000000000100010000111000000000000111110001000100000000000011100001000000001110000000011110000000001111111100000000111100001111000000000000000000000000000011010000000011111111000011101111000100000000000000000010111000000001111100000000000000001111000000000001000000000000111100000000000000000001111100001111000000001111000111110000001000000000000000000000000011110000",
		"00000000000100000000000111101110000111110000001100000000001000011111000000010000000100000001111100010000111000000000000000000000000000000000000000000001000100010001111100000000000100000000000000001111000000000000111100001111000100000000111100001111111111111111110111111110000000000000000000001110000100001110000100000000000000000000000100000000000000010000111100000001000000000000000000001111111100010001000100010000111111100000000000010001111100000000000000001111000000000000000111100000111100000000000000000000",
		"00000000000000000000000011111111000011110000000000001111000000001111000000000000000000000000000000000000000011110000000111110000000000000000000011110010000000000000000000000000000000000000000000001111000000010001111100000000000000000001000000001110111011111110111111110000000000010000000011111111000000001110000000000000111100000000000000000000111100000000000000010000000000000001000000000000111100000000000000010010111100000000111100010010000000010000000000001111111000000000000000000001111000010000000000000000",
		"11110000000000000000000000000000111111100000000000010000000100001111000000001111111100000000000000000000000000001111000000001111000100011111000000000010111100000000000011111111111100000000000000000000000011110001000000000000111100000001000000000000000011110000000000000000111100000001000000000000001000000000000000010001000000000001111100001111000000001111111100010000000011110001000000010001000011111111000000000010000011110000000000000000000100000001000000011111111111110000000000010000111100000000000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000011000001000000000000000000000000000000000000111100001111000011110000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000",
		"00000000000011111111000000000000000000000000000100000000000000000000000000100000000100001111111100000000000011111111000000000000000011110000111100000000000000000001111100000000000011110000000011100000000000000000000000000000000000000001111100000000000000011111000000000000000000010000000000010000000000010000111100000000000100000001111100001110000000010000000000000000000011110000111100000000000000000000000000000000000000001110000011100000000000010001000000000000000000000000000000000000000000000000111100000000",
		"00000000000000000000000000001111111100000001000000001111111100000000000000010000000000001111111100000000000000000000000000000000000000000001111000000000000000000000000011110000000000001111000100000000000000000001000000010000000000000000000000100001000000001111001000000000000000000000000000000001000000110000000000100000001000000010111100010000000000001111000000000000000100000000000000000000000000000000111100000001000000001111000000001111000000000000000000000001000000010000000000010010000000010000111100011111",
		"00001111000000001111000000000000111100000000000100001111000000000001000000000000000000000000000000000000000011110000000100001111000011110000000000000000000000000000000100000000000000010000111100001110000000000000000000010000111100000000111100001111000000000000000000000000111000000000000000000000000000010000111100000000000100000001000000010000000000000000000111110000001000000000000000000000000000000001000000000000000000001111000000000000000000100000111100000000000000000000111100000000000000000000111100000000",
		"00000000000111110000000000000000000000000000000100001110000000000011000000010001000000000000111100000000111100000000000000001111000000000000111100000000000000001111000100000001000000000000111100001111000111101111000000001111000011110000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000100000000000000010000000000000000000000000000001100010001000100000010000000000000111100000000000000001111000100000000000100100000000000000000000000000000111100000000000000000000111100000000",
		"11110000000100000000000100001111000000000000000100001111000000000001000000010000000000000000111100000000111000000000000000000000000000000000000000000001000000010000000011110001000000000000000000000000000111110000000000000000000000000001000000000000000000011111111100001111000000000000000000000001000000000000000000000000000000010010000000000000000000001111000000000000001000000000000000000001000000000000000000000000000000010000000100001110000100010000111100000000000011110000000000000000000000000000000000000000",
		"11110000000100000000000100000000000000000000000011111111000000000000000000010000000000000000000000000000111000000000000011110000000000000000000100000000000000001111111111110000000000000000000000000000000011010000000000000000000000000001000000000000000000010000111100010000000000001111000000000000000000000000000000000000000000000001000000000000000000001111000000001111000000000000000000000010000000000000000000000000000000000000000000001110000000010000111100000000000000000000000000000000000000010000000000001111",
		"00000000000000000001000100000000000000011111000100000000000000000000000000000000000000010000111100000001110100000000000000000000000000000001000100001111000000000000000011111111000000010001111100000000000011010000000000000000000000000000111100000000000000010001111100000000000011110000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011110001000000000000000000000000000000000000000100010000000000010000000011110000000000000000000000000000000000000000000000000000",
		"00010001000000000000000100000000000000000000000000000000000100001111000000000000000000100000000000010000110100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000011010000000011110000000011110000000000000000000000000000111100000000000111100000000000000000000011110000000000000000000000000000000000000000000000001111000000000000000000000000000100000001000000000000000000000000000000000000000000100000000000010001000011110000000000000000000000000000000000000000000000000000",
		"00000000000000000000000100000000000000000000000100000000000000000000000000000000000100010000000000000000111000000000000000000000000000010000111100000000000000000000000000000000000000000000000011110000000111010000000000000000000000000000000000000000000000000000000000000000000111110000000000010000000011100000000000000001000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000100000000000000001111111110000000000000000000000000000000000001111000011110000",
		"00010000000100000000000100000000000000000000000000000000000000000000000000000000000100010001000000100000111100010000111111110000000000010000000000000000000000000001000000000000000011110000000011100000000011100000000000000000000100000000000000000000000000010000000000000000000011110000000000000000000011100000000011111111000000000000000000000001000000000000000000000000000000000000000000000001000000010000000000000000000000001111000000000000000000000001000000000000000000000000000000010000000000000000000000000000",
		"00000000000000000000000111100000000011110000111100000000000000000000000100000000000000010001000000010000111100000000000011110000000000010000000100000001000000000010111100000001000000000000000011111111000011110000000000000000000100000000000000001111000000000000000000000000000111100000000000000001000011101111000011111111000000000000000000000001000000000000000011110001000000000001111100000001000000000000000000001101000000000000000011100000000000000001000000000000000000000000000000000001000011110000000000000000",
		"11110000001000010000000011010000111111110000110100000000000000000000000100000000000000000000000000000001000000000000000000000001000000000000000100000000000000000010000000000001000011110001000000001111000011110010000000001111000000000000000000000000000000000000000000001110000111010001000000010000000111110000000000001110000000000000000000000000111100010000000011110000000000000000111000000000000000000000000000011110000000000000000011010001000000010001000000000000000000000000000000010001000000000001000100001111",
		"00000000001000000000000011100000000000000001111000000001000000000000000100000000000000000000000011100001000011110001000000000000000100010001000000000000000000000000000000000000000011110000000000010000000100000001000011101101000000000000000000000001111100010000000000011101000111010001000000000000000000000000000000001110000000000000000000000000111100000000000000000000000000000000111100000000000011110000000000011110111000000000000011100000000000010000111100000000000000000000000000000001000000010010000100001110",
		"00000000000100010000000000010000111100000000000000000000000000000000000000010000000000001111000000000000000011100001000011111111000000010000000000000000000000001111000000000000000100000000000000010000000100000000000011111110000000000000000000000001000000000001000000010000000111100000000000011111111100000010000000000000000011110000000011011111111100000000000000010000111100000000000000000000000011110000000000001111000000000000000100000000000000000000000000000000000000000000111100000010111100000010000000001111",
		"00010000000100000000000000010001000000010000000000000000000000000001000000000000000000000000000000000000000100000000000011111111000000000000000000000000000100001111000000000000000000000000000000000000000100000000000011110000000000000000000000010000000000000000000000000010000011110001000000010000000000000010000000000000000011110000000011101111111111110000000000000000000000001111000000000000000000000000111111111111000000000000000000000000000000010000000000010000000000001111000000000011000000000010111100001101",
		"00000000000011110000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000001111000100000000000000000000000000000000000000001111000000000000000000000000000000000000000000010000000000000001000011110000000000000000000111110000000000000001000000000000000000001111000000000000000000010000000000000000000000010000000000000000000000000000000000000000111111110000000000000000111100000000000000000000000011110000000000010000000000000000000011110000000000000001000000000001000011111101",
		"00000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000100010000000000000000000100000001000000001110000000000000000000000000000011110000000000000000000011110001000000000000111100010000000000000000000100000000000000000000000000000000000000000000000000001110000000000000000000010000111111111111000000000000000000000001111111110000000011110000111000000000000000000000000000001111000000010000000000000000000000000000000000000000000000000001000000001101",
		"00000001000011100000000100000000000011110001000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000001111000000000000000000000000000000000000000000000000000011110001111100000000000000000000000000000000000000000000000100000000000000000000000000000000000000001111000000000000000000010000000011111111000000000001000000000000111100000000000000000000111000000000000000000000000000000000000000000000000000000000000011110001000000001100000000000001000000001100",
		"00000000000011100000000000000000000011100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001110000000001111111111110000000000000000111000000000000011110001000000000000111100010001000000000000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000000000000000000000000000100000000111100000000000000000000111000000000000000000000111100000000000100000000000000000000000000000001000000011100111100000000000000001011",
		"00000000000011010000000000001111000011110000000000000000000000000000000000001111000000000000000000000000000000011111000000000000000000010001000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000001111100010001000000000000000000001111000000000000000000001111000000001111000000000000000011110000000000000000000000000000000000000000000000000000111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000001100",
		"00000000000011000000000000001111000000000000111100000000000000000000000000011111111100000000000000000000111100001110111100000000000000000001000000000000000111110000000000001111000011110001000000000000000000000011000000000000111100000000000000000001000000000000000000001110000000000000111100000000000000010000000011101111000011110000000000010000000000000000000000000000000100000000111100000000111100000000111000010000000011110000000000000000000100000000000000000000000100000000111100010000000000000001000100001100",
		"00001111000011010000000000001111000011101111111000000001111100000000000100000000000000010000111111110000111100011111111000000000000011110010000000000000001000001111000000000000000000000001000011110000000011100001000011110000000000000000000000000000000000000000000000001110000000000000111100000000000100011110111111100000000000000000000000000001000000000000000000000000000000000000111000000000111100000000111100010000000011110000000000000001000000000000000000000000000100000000000000000000111100000000000000001100",
		"00000000000111100000000000000000000000000000111100010000000011111111000000000000001000100000111100001111111100000000111000001111111111100000000100000000000100010000111011110000001011110000000111110000000011110001000011101111000000001111000000011111000000010000111100000000000000000000111100001111000100011111000000000000000011110000000000000000111100000010111000000000111100000000111100000000111100000000111000010000000011110000111100100010111100000000000000000000000011101111001111110000000000000001000000001111",
		"00000000000100000000111100000000000011100000000000010000001011110000000000010000000000000000111100001111000000000000000000001110111100100001001000000001000000000000111111111111000011110000001011110000111100010001111111111111000000000000111100010000000011111111111000000000000000000001000011110000000000000000000000000000111100000001000000000000111100010000111100100000110100000000000100000000000000000000000000000000000100001111000000000001111100000000000000001110111111100000000011100000111000000001111100010000",
		"11100000000000010000000000001111000000000000111100010000000000001111000000001111000000000000111100000000000011100000000111110000000000100000000011110010000000000000000000000000000011110000000111111111111100000001111100000000000000000001111100001110111011111111111100000000111100000000000000000000000000001111111100000001000000010000000011110000111100010000111100000000000000000000000000000001111000000000000000010010000000000000000100000000000100011111000000001111111100000000000000000001111100010000000000000000",
		"11100000000000100000000000010000000000000000000000001111000011111111000011111111111100000000111100000001000000001111001000000000000100011111111100000001000000000000111100000000000000001111111111110000000000010001000000000000111100010001000000010000000011101111000000010000000000000001111100000000000100010000000000000010000000010010111100001111000000000000000000000000000111110001000000000001111100000000000000000001000011110000000111110000000100000000000000001111000000000000000000000000111000000000000000000000",
		"00000000000000000000000000010000000000000000000000000000000011100000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001111000000000000000011110000111100000000000000000000000000000000000000000000000011110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
		"00100000000000000000000000001111000000000000000000000001000000001111000000001111000000000000000000001111001000010000000000010000000000000000001011101111000100010001000000000001000000000000000011100000000000000000000000000000000000000000000000000000000100011111001011100000000000011111111100010000000100000001000011110000000000001111111100011110000100000000000000010000000000010000111100000000000000000000000000001111111111110000111111111111000000000001000000000000000000000000000000000000001000010000000011110000",
		"00000000000000000000000000001111111000000001111100000001000011110000111100010000000100000000000100100001000000001111000000000000000000011111000000000001000000000000000000001110111100001111000011110001111100000001000000000001111100000000000000000001000000000000000000001111000000000000000000000000000000000001111111110000000000000001111100000000000000000001111011100000111100000001000011110000000100000000000011110000111100000000000000000000000000100001000000011111000011110000000000100000111100000001000100000000",
		"00000000111100100000000000001111000000000000000000001111000000000001000000010000000000000000000000000001000000001111000011110000000000010000111100000000000000011111001000000000111100000000000000000000000000000001000000000000111100000001111100100000000000010000000000000000000000000000111111110000000000010000000000010000000000000001111100000000000000001111000000000000000111110000000000000000000000000000111100000000111100001110000011111110001000100000000000000000000100100001111100010010000000000000000011111111",
		"00001111000100001111000011110000000000001111000000001111000000000010000100000001000000000000000011110001111111110000000100000000000000000000111100000000000000001111001000000000000000000000000000001110000000000001000000000000111111110000000000001110000000000000111100010000111100000000000011110000111100010000000000000000000000010000111100000001111100000000000000000000000000000000000100000000000000000001000000000000111000001111000100000000001000010000000000000000000000000000111100000000000000000000111100000000",
		"00000000000100000001000011111111000000000000000011111111000000000001000000000001001000000001000000000000111100000000000100000000000100000000111000000000000000011111000000000000000000000000111100001110000011010000111100000000000011100000000000000000000000000000111000010000111111110000000000000000000000000000111100011111000000000001000000000001000000000000000100000000001000010001001000000001000000000000000000000000111100000000001000000000000100000000000000010000000000000000000000010000000000000000000000000000",
		"00000000000000000000000100000000000000000000000111111111111100000001000000010000000100100000000000100000111100000000000000000000000000000000111100000000111100000000111100000001000011110000000000001111000111010000000000000000000011110001000000000000000000001111111100000000000000001111000000000000000000000000000000010000000000010010000100000000000011110000000000000000000100000001000111110000000000001111000000000000000000000000000100001110000000001111000000000000000011110000000100000000000100000000000000000000",
		"00000000000000000001000011110000000000000000000011100001000000000000000000011111111100100000000000000000111100000000000000000000000000000000000100000000000000000000000000000000000000000000111100000000000011000001000000000000000011110000111100000000000000010000000000000000000000000000000000000000000111110000000000001111000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000111100000000000000001111000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000000001000011100000000000000000000011110000000100000000111100000000000000010000000000000000111000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000011000000000011110000000100000001111000010000000000010000000000010001000011110000000000000000000011100000000000000000000000000000000100000000000000001111000000000000000011110001000100000001000000001111000000000000111100000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000",
		"00000000000000000000001011100000000000000001000111110000000000000000000000000000000100100001000000000000111100000000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000111100000000011110000000000000000111100010000000000000000000000010000000111110000000000000000000011110000111100000000000000000000000100000000000000000000000000000000000000000000000100000001000100000000000000000000111000000001000100100000000000000001111100000000000000000000111100000000000000001111000000000000",
		"00010001000000000000000111100000000000000000000000000001000000000000000000010000000100010000000000010000000000100000000000000000000000000000000000000000111100000001000000000000000000000000000000000000000011110000000011110000000000000000000000000000000000000000000000000000000011110000000000000000000011100000000011110000000100000000000000000001000000000000000000000000000000000000000100000000000000010000000000001111111100000000000100010000000000000001000000000000000011110000111100000000000011111101000000001111",
		"00000001000000000000000111100000000011110001000011110000000000000000000000000000000100000001000000010001000000000000000000000000000000011111000000000001000000000001000000000000000011110000000011110000000100000000111100000000000000000000000000000000000000010000000000000000000111110000000000000000000011110000000011101111000000000000000000000010000000010000000000000000000000000000000000000001000000000000000000001111111111110000000000010000000000000001000000001111000000000000000000010001000011101111000000000000",
		"00000001000000000000000011100001000011110000111000000000000000000000000000000001000000010010000011110001000100000000000011111111000000000000000000000001000000000001000011110001000000000001000000000000000000000000000000000000000100000000000000001111000000000000000100000000000111110000000100000000000000000000000000001101000000000000000000000001111100000000111111100001000000000000000000000000000000000000000000001101111111110000000000000000000000010001000000000000000000000000000000010000000011100000000000010000",
		"00000000000100000000000011010001000000000001111000000000000000000000000000000000111100000000000011110001000111110000000000000000000000010000000000000001000000000001000000000000000011110001000000010000000000000001000000001111000000000000000000000000000000010000000100001111000111110001000000001110000000010000000000011110000000000000000000000000000000000000111100000001111100000000111100001110000000000000000000001101110111110000111111110001000000000001000000001111111100000000000000000000111100000010000000000000",
		"00000000000000000000000000000000000000000001111100000000000000000000000011110000111100001101000011100000000011110001000111111111000100000000000000000000000100001111000100000000000011100000000000000000000100000000000011111110000000000000000000000000000000010000000000001111000011110000000011111110000000010000000000000000000000000000111011110000111111110000000000010000111100000000000000001110000000000000111100011111110100000000000000000000000000000000111000000000000000000000000000010001111100100001000100000000",
		"00000000000100000000000000010000000000000000000000000000000000000000000000000000111100001111000000000000000011110001000011110000000100000000000000000000000000001111000100000000000000000000000000000000000100000001000000000000111100000000000000000000000011110000111100010000000000000000111100001111111000000001111100010000000000000000111011010000111011110000000000000000111100001111000000001111000000000000000000001111111100000000000100000000000000000000111100000000000000000000000000000001111100000001000000000000",
		"00000000000000001111000100010001000000000001000011110000000000000000000000000000111100100000000000000000000000000000000011110000000000000000000000000000000000001111000100000000000000000000000000000000000000000001000011110000000011110000000000000000000011110000000000010010000000000000000011110000111100000001000000000000000011110000111111100000111100000000000000000000111100001111000000001111000000000000000011110000000000000000000000000000000000000000111100000000000000000000000000000001000011110010000000000000",
		"00000000000000000000000100000001000000000000000000000001000000000000000000000000111100010000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000010000111100000000000000000000000000000000000011110000000000000001000000010000000111110000111100010000000000000000000000000000000000001111000011110000000011110000111011110000000000001111000011110000000000000000000000000000000000000000000011110000000000000010111111110000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000011110001000000000000000000001111000000000001000000010000000000000000000100000001000000000000000000000000000000000000110100000000000000000000000011110000000100010001000000000000000000000000000011111110000000000001000011110000",
		"00000000000011110000000000000000000000000001000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100001111000011110000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000001000000000000000000001110000000000000111100000000000000000000000000000000000100000000000000000000000000000000111000000000000000000000000000001111000100000001000100000000000000000000000000001101000000000001000011111110",
		"00000000000011100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010001000111110000000000000000000000001110000000001111111100000000000000000000111100000000000011100000111100000001000000100001000000000000000000001111000000000001111100000000000000000000111100000000000000000000111100000000000011110001000100000000000100000000000000000000000011110000110100000000000000010000111100000000000000000000000000000000000000000000111100001110111100000000000000001110",
		"00000000000011010000000000000000000000000001111100001111000000001111000000000000000000010000000011110000000000000000111100010000000100000000001000000000000011111110000000000000000000001111000000000000111111110000000011110000000000000000000000100000000000000000000000011111000000000001111100000000000000000000000000010000000000000000111100000000000000000001000100000000000000000000000000000000000000000000110100000000000000010000111100000000000100000000000000000000000011111110000000001110000000000000000000001101",
		"00000000000011010000000000001111000000000000000000000000000000001111000000010000000000010000000000000000000100001111000000010000000000000001000100000000000000001101000000001111000000000000000000000001111111110010000000000000111100000000000000010000000011110000000000001110000100000000111000000000000000001111000000000000000011110000000000000000000000000000000100000001000000000000000000000000111100000000110000000001000000000001111000000001000011110000000000000000000000001111000000001111111100000000000000001100",
		"00000000000011000000000000011111000000000000111100100000000000000000000000001111000100010000111100001111000000001110000000000001000011110010000000000000000000001110111100001110000000000000000000000000111111110001000011110000000000000000000000000000000000000000000000001110000000000000111000000000000000000000111100000000000000000000111100000000111100000001111100000000000000100000000000000000111100001111110100100001000000000000111100000011000011100000000000000000000011111110000000000000000000000001000000001101",
		"00001111000011010000000000011110000100001111111100101110000000001111000011101111010000100000111011110000110100010000111100000000000011110010000000000000000100000000111100000000001011110001000011110001111100000001000011111111000000000000111100010000000100010000111100001111000000000000111100001111001000001111111000101111000011101111000000000001000011110010111000000000111100100000000011110000111000011111110100100001000000000000111100000010111111100000000011111111000011111101001111110000000000000010000000001110",
		"00001111000011110000000000001111000111100000111000111110000000000000000000000000001000001110111011110000110100000001000000000000000000010001000011110000000100001111111100000000000011110000000000000000000000000000111111101111000000000001111000001111000000001111111111110000000000001111000011110001000111110000111100001111111100010000000100000001000000000001111100000000111000010000000011110000110100000000000000010000000100101111000000000000000000000000111100001111000000001111000111110000000000010000000000001111",
		"00001111000000010000000111111110000000000000111100000000111100001111000100000000000100000000111011110001111100000000000111110000000100000000111100000010001000000000000000000000001011100000000000000000000000000010111100000000000000000001111000000000000000000001111111110000000100001111000000000000000000001110111000001111000000010000000000000001000000000000000011100000000000000001000011101111111000000000000000010001111111110000000000000000000100001110000000001111000100010000000000000010111100100010000111100000",
		"00001111000000100000000000011111000000010000000011110000000100000000000011111110111100000000111100000001000100010000000100000000000100000000000000000001000000000000111100000000000011110000000011100000111100010001000000000000111000000001111100010000000000001111000000000000000011110010111111111111000000010000000000010001000000100001111100000000111100000001000000000000000000000000000000000000111100000000000000000000111111111110000111111111000100000000000000001110000100000000000011110000111000100001000000000000",
		"00000000000000001111000000010000111100000001000000000000000011110000111100000000111100000001000100000000000000001111000000000000000000010000000100000001111100000000111111110000111111111111111111100001111100000001000000000001111100000010000000000000111000000000111100001111111100000001000000011111000100000001111111110001111100000000111100011111000100010000111100010000000011110000000000000000000100001111000111100001000100000001000011111111000100000001111100011111000011110000111100010000111100010000111100000000",
		"00000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000001000100000000000000000000111100000000000000000001000011110001000000010000000100000000000000010000000000001110000000010000000000001111111100000010000000000000000111111111000000000000000000000001000000000001000000000000111100000001111100000000000000000000000000000000111100000000000000000000000000000001111100000000000000000001111100000000000000010000000011110000111100000000000000000000000000001111000000000000000000001111000100001111000000100000000000011111000011110000000000010000111100000001000000000000",
		"00010000111100001111001000000000000000100000001000000000000011110001000000100000000000010000111100000000111100000000000011111110000100000000000000000000000100011111000100010001000000000001000000000000000100000000000011111111000011110010111100001111000000001111111100010000000000000000111011110000111100000000000000000000000000000010000000010000000000001111000011111111000000000000000100001111000000000000000000000000111000001111000000000000000100100000111100010000000000000000000000010000000011110000000011100000",
		"00000000000000000000000011101111000000001111000011110000111100000001000100000000000000000000000000000000111100000000000000000000000000000000111000000001000000010000000000000000111100000000111100000000000111100001000100000000000000000001000000000000000000000000111100010000111111110000111100000000111100010000000000000000000000000001111100000010111100000001000100001111000000000000000100000000111100000000000000001111110100011110000011110000001100000000000000000000000000000000111100100000000000000000111100000000",
		"00000000000000000000000011101110000100000000000011110000111100010010000000000001000100010001111100000000000000000000000011110000001000000000111100000000000000000000000000000000000000000000000000000000000111010000000000000000000011110010000000001111000000000000000000000000000011100000000000000001111100000000000000001111000000000010000100000000000000000000000000000000001000010000000100000000000000000000000000011111110100000000001000000000000100000000000000010000000000000000000000010000000000000000000011110000",
		"00000000000000000000000111101111000100000000000111111111111000000000000000000000000100110001000000010000000000000000000000000000000000000000111100000000000000000000111100000000000000000000000000000000000011010000000000000000000000000001000011110000000000010000000000010000000011110000000000000000000000000000000000001111000000000001000100000000111100000000000011110000000100010001000100000000000000000000000000001111110100000000000100000000000000000000000000000000000000000000000000001111000011110000000011110000",
		"00000000000000000000000011011111000000000000000011110000000000000000000000000000000000100000000000000000000000000000000000000000000000010001000000000000000000000000000011110000000000000000000000000000000011110000000000000000000000000001111100010000000000000000000000010000000111110000000000001111000011100000000000001110000000000001000100000000000000000000000000000000000000000001000100000000000000001111000000001111110100000000000000010000000000000001000000000000000000000000000000000000000011110000000000000000",
		"00000000000011110000000111000000000000000000000000000000000011110000000000000000000000010001000000000000000000011111000000000000000000000000000000000001000000000000000000000000000000000000000000000000000011110000000000000000000011110001111100010000000000000000000000100000000000000000000000001111000011100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000110100000000000000011111000000000001000000000000000011110000000000000000000011110000000000010000",
		"00000000000000000000000111000000000000000000000011110000000000000000000000000000000100010000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000011110000000100001111000000001111000000000000000000000000000000000000000100010000000100000000000000000000000011110000000000001111000000000000000100000000000000000000000000000000000000000001000100000000000100000000000000001111110100000000000100010001000000000001000000000000000000000000000000000000000000001111000000000000",
		"00000000000000000000000011010000000000000001000000000000000000000001000000000000000000000001000000000000001000000000000000000000000000010000000000000000000000000001000011110000000100000000000011110000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000001110000100000000000100000001000000000000000000000000000000000000000100011111000100000000000000001111111000000000000000100000000000000001000000000000000000000000000000000000000000001110000000000000",
		"00000000000000001111000011100001000000000000111100010000000000000000000000000000000000000010000100000000001011100000111100000000000000000000000000000000000000000001000000000000000000000000000011100000000000010000000000000000000100001111000000001111000000000001000000010000000000000000000000000000000000000000000000001111000011110000000000000010000000010000000011110001000000000000000100011110000100010000000000001110111011110000111100010000000000000001111100000000000000000000000000000000000011111111000000000000",
		"00000000111100011111111111110001000000000000111000010000000000000000000000000000111100000010000011110000001011100000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000010001000000000000000000001111000100001111000000000000000100000000000111110000000100001110000000010000000000001111000000001111000000000000000000010000111000000001000000010000000000011101000100000000000000001110111011100001000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
		"00000000111000001111000000000001000000000000111100010000111111110000111111110000111000000000000011110000000011100000000000000000000000000000000000000000000100000000000000000000000100000000000000010000000000010001000000000000000011111111001000000000000000000000000000000000000100000000000111111101111100010000000100011110000000000000000000000000000000001111111100000001000000000000111100011101000000000000000000001110111000000000111011110001000100001111000000000000000100010000000100000000000000010000000000000000",
		"11110000111000000000000000000000000000000000111100000000000011110000111100000000111000001101000000000000000011110010000011110000000000000001000000000001000000001111000100000000111111110000000000000000000000000000000000000000111111110000000100000000000000000000000000000000000000000001000011110000111000000000000000000000000000000000000011100000111100000000000000100001111100000000000000001111000000000000111100000000111100000000000011110000000011110000000000000001111100000000000000000001111100010001000000000000",
		"00000001111100000000000100000001000000000001000000000000000011110000000000000000111000010000000000000000000000000001000011100000000100000000000000000001000000001111000100001111000000000000000000000000000100000001000000000000000011100000000000000000111111110000111000000000000000000001000000000001111100000001000000000000000000000000111111000000000000000000000000010000000011111111000000000000000000000000000011110000000000000000000000000001000000000001000000000001000000000001000000000000111000000001000000000000",
		"00000000000000001110000100000010000000000001000000000000000000000000111100000001111100000000000000000000000000000000000011010000000000000000000000000000000000001111000000000000111100011111000000010000000000000000000000000001111111110000000100001111111000000001111100000000111100000000000100000000111100000001000000000001000011110000111111100000000000000000000000010000000000000000000000000000000000001111000011100000000000001111000000000000000000000001000000000000000000000000000011110000000011110001000000000000",
		"00000000000000000000000000000001000000000000000000000000111100000000000000000000111100000000000000000000000000000000000111110000000000000000000000000000000000000000000100000000111100010000000000000000000000000000000000000001000000000000000000010000111100000000000000000000000000000000000011110001000000000001000000001111000011110000111100010000000000000000000000000000000100000000000000000000000000000000000011110000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000111110000",
		"00000000000000000000000000000001000000000000000000000000000000000001000000010000000000000000000000000001000000000000000011110000000100000000000000000000111100000000000000000000000000001111000000000000000000000000000000000000111100000000000000000001000000000000000000000000000000000000000000000001000000000001000000001110000000000001000000010000000000000000000000000000000100000000000000000000000000000000000000000000111100001111000011111110000100000001000100000000000000000000000000001111000000000000000011110000",
		"00000000111100000001000000000001000000000000000011110000000000000000000100010000000000000000000000000000000000000000000000000000000100001111000000000000111100001110000000000000000000001111000000000001000000000000000000000000000011110000111100010001000100000000000000001111000000000000000000000001000000000000111100001111000000000000111100000001000000000000000000000000000100000000000000010000000100000000111000000000111100000000000000001110000000000000000000000000000000000001000000001110000000000001000011110000",
		"00000000111100000001000000000000000000000001000000000000111111110000000000000000000000010000000000000000000000000000000000000000000000001111000000000000000011111111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000000000000000000000000000000000001111000000000000000000000000000011110000000000000000000111110000000000010000000000000000111000000000000000010001000000000000000000000001000000000000000000000000000000001111000000000000000011110000",
		"00001111000011110001000000000000000000010010000000001111000011111111000000000000000000010000000000000000000100000000000000000000000100000000000100000000111111111111111100000000000000001111000000000000111000000000000000000000000011110001000000000000000100000000000000000000000100000000000000000000000011111111000000000000000100000000000000000000000000000001000100010000000000000000000000000000000000000000110100000000000000010001000000000000000100000000111100000000000011111111000000001111000000000000000000000000",
		"00000000000011100000000000000000000000000001000000000000111100000000000000000000000100000000000000000000001000001111000000000000000000000001000100000000111100001111111100001111000000001111000000000000000011110000000000010000000011100000000000000000000000001111000000001111000000001111000000010000000011111111000011111111000000001111111100000000000011110000000100000000001000000000000000000000000000000000111000000000111100000001111100000000000011110000111100000000000011111110000000011111000000000000000000001111",
		"00000000111111100000000000000000000000000000000000010000000000000000000000001111001000001111000000010000000000001111000000000010000100000010000000000000000000001111111000001111000000000000111100000000000011110001000100000000000011110001000000000000000000010000000000011111000000000000111000000000000000001111000000000000111100000000111000000000000011100001000011110000001000010000000011111110111100011111111000010000111100010001111100010010000011100000111100000000000000001110000000000000000111110010000111101111",
		"00001111000011010000000000011111000100011111111100011100000000001111000000001111000111110000111100000000111100010000000000000000000000000001000000000000001100001111111100000000000100000000000000000000000000000000000011100001000000000001000000001110001000011110000000010000000000001111111100000000000000001111111000000000000011111111110100000000000011100000111100001110000100100001000000001111111100001111111000000001000000000000111100000001111111100000000000010001000111111110001000000010000100010000000011111111",
		"00100000000011111111000000011110000000001111111100011101001000000000000000001111000011111111111011100000111100001111000000000000000000100000000100000000001000001111000000000000000000000001000100001110111100100000111111110000000000000001111000001110000000001101111100000000111111110000000011101111000000011110111111110000111100011111111100000000111111110000110100010000000000010000000000000000111000000000000000000001000000011110000000000000000000000000111100001111111111101111000011110001000000100000000000101110",
		"00000000000100000000000000001110111111110000000000100000000011110000000100001111000011110000111000000000000011101111000011110000000000100001000111100010000100000000000000000000000011010000001011111111111100100000111000000001111100000010111000001110111000001110111100000001111100000000000000001111000000000000000000010000000000010001000011111111110100000000111100000000111100011111111100000000111000000000111100000000000000001101000100000000000000000001000000001101111111110000000000000000111000010001000000000000",
		"00001111000000011111000000001110000011110000000000000000001000000000000011111110111011110000000000000001000100001111001000000000000100010000000000000010000000000000000000001111111011100000000011110000111111100000000000000000111000000001111000000000000000101111000000000000111000000010111100001110000000010000000000000000000000010001111100001111111100001111111100101111111111110000000000100000111011110000000011110000000000001110000011101111001000000001000000011110111111101111111100000001111000110000000000010000",
		"11111111000100010000000000001111000100010000111100001111000000001111000011110000000011110000000000000000000011110000000000000001000000000000000000000000000011110001111100011111000100010000000000001111000000000000111100000000000000010000000111110000000000000001000000010000000111110001000000001111111100000000111111110001111100010000000000000000000000000000000000001111000000000000000000011111111100000000000011111111000000000000000000000001111100000000111100000000000000000000000011110000000000010001111111110000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000",
		"00000000000000001111000000001111111100000000000000010000000000000001000000010000000000000000000000000000000100001110000000000000000000010000000011110000000000000000000000001111111111110000111111100000111100000001000000000000111100000000000000000000000000000000000011110000111100000000000000001110000000000000000000000001000000000000000000000000000000010000111100000000000000000000000000000000000000000000000000000000000011111111000000001111000000010001000000010000000011110000000000000001111100010001000000000000",
		"00100000000000010000000111111111000100000000000000001110000011110000000100010000000000000000000000000001000000000000000011111110000100000000111100000000000000000000000100010000000011110001000100000000000100000000000000001111000000000001000000000000000000010000111100010000000000000000000011111111111100000001000000010000000000010010000000000000111100001111111100001110000000001111000000011110111111110000000000001111111000000000000011110000001000010000000000011111000000010000000000100000111100000000111111110000",
		"00000000111100000000000011001111000000000000000011111111000000000001000000010000000000000000000000100001111100010000000000000000000100000000110100000000000000010000000000000000000011110000111100000000000011110001000100000000000000000001000011110000000000000000000000010000000000000001111100000000111000000000000011100000000000000010000000000000000000000000000000001111000000001111000100001110111100000000000000001101110100001110000011111111001000000001000000010000000000001111000000100000111111110000111000000000",
		"00000000000011110000000111011111000000000001000000000000111000000001000000000001000000100001000000000000000000001111000011110000000100000000000000000000000000000000111100000000000000000000000000000000000011110000000000000000000011110010000000000000111100001110000000100000000000000000000000000000111100000000000011111111000000000010000000000001000000000000000000000000000000000000000100001111000000000000000000001110110000000000000000001110000111110000000000010000000000000000000000011111000000000000111100000000",
		"00000000000000000000000011010000000000000000000000000000111100000000000000000000000000010001000000000000000000001111000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000010111100000000000000000000000000010001000011110000000000000000000011100000000000001101000000000001000000000000000000000000000000000000000100000001000000000000000000000000000000001111110000000000000000001111000011110001000000010000000000001111000000010000000011110001000011110000",
		"00000001000000000000000011000000000000000000000000000000000011110000000000000000001000000000000000000000000000000000111100000000000000010000000000000001000000000000000000000000000000000000000011110000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000111111110001000100001110000011110001000100000000000000000000000011110000000000000000000100001111000000000000000000001111110000000000111100010000111100000000111100000000000000000000000000000000000011110000000000000000",
		"00000000111100000000000011100000000000000000000000000000000000000000000000000000000100000001000000000000000000010000111100000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000011110000000000000000000000010000000000000000000000000000000100000000000000001111000000000000000000001110000000000000000100000000000000000000000000000000000000000000000000000000000100001111000000000000110100000000000000000000111111110001111100000000000000000000000011110000000011110000000000000000",
		"00000000000000000000000011100001000000000000000000000000000000000000000000000000000100000001000000000000000100000000000000000000111100000000000100000000000100000001000000000000000100000000000000000000000000010000000000001111000000000000000000000000000000000000000000000000000100000000000000001111000000000000000000001110000000000000000100000000000000000000000011110001000000010000000000001111000100000000000000000000111000000000000000010001000000000001111100000000000000000000000000000000000011110000000100000000",
		"00000001000000000000000011110010000000000000000000010000000000000000000000000000000100000001000000001111001000000000111100000000000000000000000000001111000000000000111100000000000000010000000011110000000000100000000000000000000000001111000000000000000000000000000000000000000000000000000100000000000000000000000000001111000011110000000000010000000000000000111111110001000000001111000000001101000100010000000000000000111100000000000000010000000000000000000000000000000100000000000000010000000011111111000000000000",
		"00000000111100000000111100000001000000000000111100010000000000000000000000000000000100000010000011110000000111100000000000000000000000000000000000001111000000000000000000000000000000000000000111110000000000010001000000000000000100001111000000000000111100000000000000000000000000000000000100000000000000010000000000001111000011111111000000010001000100000000000000000001000000000000000000001100000000011111000000000000111100000001111100010000000000000000000000000000000100000001000100010000000011110000000000010000",
		"11110000111000000000000000000000000000000000111000000000111100000000111111110000000011110000000011110000000011100000000000000000000000000000000000001111000011110000000011110000000000000000000000000000000000010001000000000000000000001111000100000000000000000000000000000000000000000000000100000000111100010000000100000000000011111111000100010000000000000000111000000000111100010000000000001101000000001111000000000000000000000000111000000000000000001111000000000000000100000000000100000000000100000000000100100000",
		"00000000110000000000000000000000000000000000111100000000111100000000111111110000000000001110111100000000000000000001000000000000000000000001000000000000000011111111000000000000000000000000000000000000000000000000111100001111000100001111000100000000000000000000000000000000000000000000000000000000111100001111000100000000000100010000000100000000000011110000000000100001111100000000000000000000000000000000111100000000000000000000111000000000000011111110000000000001000000010000000000000000000100010000000000010000",
		"00000000111100000000000000000000000000000000111000000000000011110000000011110001000000001101111100000000000000000001000100000001000000000001000000000001000000001111000000000000000000000000111100000000000000000000111100000000000011111111000100000000000011110000111100000000000000010000000100000001111100000000000000000000000000100000000011100000000011110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000000001000000000000000000000000000000000000",
		"00000000111100001111000100000001000000000001000011110000000000000000000000000000000000000000000111110000000000010000000011110000000000000000000000000001111111110000000000000000000000000000000000010000000000000000000000000000000011110000000000001111111100000001111000000000000000000000000100000001000000000000000000000000000000000000000011000000000100000000000000000000000011111111000000000000000000000000000100000000000000000001000000000001000000000000000000000000000000010000000000000000000000000000000000000000",
		"00000000000000001110000000000010000000000001000011110000000000000000111111110001000000010000000000000000000000000000000011100000000100001111000000000000111100000000000000001111000000010000000000010000000000000000000000000000000000000000000100000000111100000001000000000000000011110000000000000000111100000000000000000000111100000000000000000000000000000000000000010001000100000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000",
		"00000000000000000000000000000001000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011100000000100000000000000000000000011110000000000000000000000010000000000000000000000000000000000000000000000000000000000010000111000000001000000000000111100000000000100000000111100000001000000000000000000000000000000010000000000000000000000000001000100000000000000000000000011110000000011110000000000001111000000000000000000010000000000000000000000000000000011110000000000000000000000000000",
		"00000001000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000100000000000000000000000011111111000000000000000000010000000000000000000100000000000000000000000000000001000000010000000000000001000000000000111100000000000100000000111100000001000011110000000000000000000000000000000100000000000000000001000100000000000100010000000000000000000000000000111100000000000000001111000100000000000100000001000100000000000000000000000000000000000000000000",
		"00010000111100000001000000000001000000000000000011110000000000000000000000000000000000000000000000000000000000000000111100001111000100000000111100000000000000000000000000000000000000001111000000000001000000000000000000000000000000000000000000000001000000010000000000000000111100000000000000000000000000000000000000001111000000000000000000000001000000000000000100010000000000000000000100011111000100000000000000000000000000000000000000001111000000000000000000000001000000000001111100001110000000000000000011110000",
		"00000000111100010001000100000001000000000001000011100000000011111111000000000000000000010000000000000000000000000000000000001111000100001111000000000001000011101111000000000000000000001111111100000000000000000000000000000000000000000000111100010000000000000000111000000000000000000000000100000000000000000000000000000000111111111111000000000000000000000000000000010000000011111110000100010000000000000000000000001111000000010001000000000000000000000000000000000000111100000000000000001110000000000000000011110000",
		"00001111000000000000000100000000000000000010000011110000000000001111000000000000000000010000000000000000000000001111000000011111000000000000111100000000111000000000111100000000000000001111000000000000111100001111000000000000000011110001000000010000000000001111111100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000100000000000000001111000000000000000000000000000000000000000000010000000000010000000000000000000000010000000011111111000000000000000000000000000000000000",
		"00001111000011110001000000001111000000010001000100000000111000000000000000000000000100100000000000000000000000001111000000001111000011100000000000000000111111110000111100000000000000001111111100000000000000000000000000010000000111110010000000000000000000000000000000000001000000001111000000010000000011100000000111110000000000001111111100000000000000000000000100000000001000010000000000000000000000010000000000000000000000100000111100010000000000000000000000000000000111101111000000010000001011100000000011110000",
		"00000000000000000000000000001110000000010000000000011111000000010000111100000000000100010000000000000001000000010000000000000000000011110001000000000000000011110000111100000000000000000000111100001111000000000000000000001111000111110010000011110000000100011111000000000001111111110000000000000001000011101111000011110000000000001110111100000000000111110000000000000000001000100000000000010000000000101111111000000000000000010000111100000000000011100000000000000001000011111111000000010000001011110000000011110000",
		"00000000000000001110000000011111000000000000000000011101000000000000000000001111000000000000111100000001000000010000000000000000000000010000000000000001001000010000111100000000000000000000000000000000000000010000000000000000000000000010111100000000000000011101000000100000111111111111000000000000000011110001000011100001000000001111111000000000111111110000110100011111000100100000000000010000000000001110111100000000000000011111111100000000111111100001000000100000000011101111000000010001000100001111000000000000",
		"00000000000011111111000000000000000000011111000000001110000000000000000000001111000011101111111100000000000000011111000100000000000100010000000100000001000100010000111100000000000000000001000100001111000000100000000000000001111100000001110100001111000000001110111100000000000011110000000011111111111100000000111111110000000000001111111100000000000011111111110100000000000000000000111100000000000000001111111100000000000000001111111100000000000000000000000000100000000011101111000000010011000000010000000000001111",
		"11110000000000000001111100001111000011111111000000010000000000000001000000000000000011110000111100001110000000000000000011110000000100011111000111100000000100000000000000000001000011100000001000011111111100010000111100000001000000010010111000001111000000001110111100000000111100001111000111110000000000000001000000000000000000000000000011111111110100001111111100000001000000010000111100000000000011110000111100000000000000101110000011111111000000000000000000011111000011110000000000000001000000010000000000011111",
		"00000000000000000000000000000000000000000000000000000000000000010000000000000000000011110000111100000000000000000000000000000000000000011111000000000000000100000000000000000000000000000000000100000000000000000000111111110000000000000000000000000000000100000000000000000000111100000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000010000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000100000000000000000000111100000000111100000000000011110000000100000000000000000000000000000000000100001111000000000000000000000000111100000000000000000001000000010000000000001111000011110001111100000000000000000001000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001000000010000000000000000000000000000111100000000000000000000111100000000000000000001000000000000000011110000000100000000000000010001000000000000000000000000000000000000000000000001000000000000",
		"00010000000100010000000000001111000000000000000000001110000000000000000000000000000000000000000000000000000100000000111100000000000000010000111100000000000000000000000000011111111100000000001000000000000100010000000000000000000000000000000000000000000100000000111100010000000000000001000011111111111000000000111100010000000000010001000000001111111100001101000000010000000011110000000000011110000000000000000000000000111000000000000011110000000100000001000000011111000000010000111100000000000000000000111100000000",
		"11110001111100000000000011101111000000000000000111110000000000000001000000000001000100000000000000110000000000011110111100000000000000010000111100000001000100000001000000001111000011110000000000000000111100010000000000000000000000000001000000000000000111111111111100010000000000000001000011110000111100000001000011111111111100000010000000000001000000001111000000010001000011110000000100001111000000000000000011111110111100001111111100001111000100001111000000000000000011100000000000000000000000000010000000010001",
		"00000000000011110000000011111111000000000000000000000000111100000001000000000000000000010001000000010000000000001110000000000000000000000000000000000000111100000001111000000000000000001111000000000000111100000000000000000000000000010010000000000000000000001111000000010000000000000000000000001111000011110000111111101110111111100000000000000000000000000000000000000000000000010000000000001110000000000000000000011110111000000000110100001111000011110001000000000000000011110000000000001111000011110001000000000000",
		"00010000000000000000111100000000000000000000000100001111000000000000000000000000000000010000111100000000000000000000111100000000000000000000000000000000000000010000000000000001000000001111000000000000000000010000000000000000000000000010111100010000000100000000000000010001000000000000000011110000111111110000000000001101000000000001000000000000000000000000000000000000000000010000000000001110000000000000000000010000111000000000111000001111111111110000000000000000000000000000000000001111000000000010000000000000",
		"00000001000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001000011110000000000001111000100000000000000011111000000000000000000000001000000000000000000000000000000000001000100000000000000000000000011100000000000001110000011110000000000000000000100000000000000000001000000000001000100001110000000000000000000000000111000000000111100000000000011110000111100000000000000000000000000000000000011110000000000000000",
		"00000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000010000111100000000000000000000000000001111000000000001000000000000000000001111000100000000111100100000000000000000000000000001000000010000000000000000000000000001000100000000000000001111111000001111000000001111111111110000000000000000000000000000111100000001000000001111000000011111000000001111000000000000111100000000110100000000111111110000111000000000000000000000000000000000000011110000000000000000",
		"00000000000000000000111100000001000000000000000000010000000011110000000000000000000000000001001000000000000100000000000000000000111100000000000000001111000000000000000011110000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000001000000000000000000000000111100000000000000000000000011110000000000000001000000000001000000000001000000001110000000001110000000010000000000000000000100010000110100000000000011100000111100000000000000001111000100000000000011110000000100010000",
		"00000000000000000000000000000001000000000000000000100000000000000000000000001111000100000001000100000000000111110000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100010000000000000000000000000000000100000000111100010000000000000000000000001111000000000000000000000000000000000000000011110000000100000000000000000000000000000001000000001110000100001110000000011111000000000000000000000000111000000000000011100000000000000000000100000000000000000000000000000000000000010000",
		"11110000111111100000000000010000000011110000000000010000000000000000111111110000000000000000000011110000000011100000000000000000000000000000000000001111000000001111000000000000000000010000000011110000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000011101111000000010001000100000000000000000000000000000000000000000000000000010000000000000000000000000000111000010000000011110000111100000000000000000000000100000000000000000000000000010000",
		"00000000110100000000000000010000000000000000111100000000000000000000000000000001000000001110000000000000000000000000000000000000000000000001000000001111000011110000000011110000000000010000000000000000000000000000000000000000000000001111000100000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000100000000000000100001000000001111000000000000000000000000000000000001000100000000111000000000000011111111000011110000000000000001000000000000000000010000000000100000",
		"00000000111000000000000000000000000000000001111100000000000000000000000000000000000111111101000000001111000000000000000100000000000000000000000000000000000011110000000000000000000000000000000000011111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000011110001000000001111000000000000000000010000000000000000000111110000000000010001000011110000000000000000000000000001000000000001000000000000111000000001000000001111000000000000000000000001000000000000000000100000000000010000",
		"00000000111100010000000000000000000000000000111000000000000100000000000000000000000000001110000000000000000000000001000000000000000000000000000000000001111111111111000000000000000000000000111100010000000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000000011111000000000000000000010000000111100000000100000000000000000000000011111111000000000000111100000000000000000000000000000001000000000000000000000000000011110000000000010001000000000000000000010000000000000000",
		"00000000000000001111000100000000000000000000111100000000000000000000000011110000000000000000000000000000000000010000000000000000000000010000000000000000000011110000000000000000000000010000000000000000000000000000000000000000000011110000000000000000000000000000111100000000000000000000000100000000000000000000000000000000111100000000000011010000000100000000000000000000000100001111000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010001000000000000000000000000000100010000",
		"00000000000000000000000100000001000000000000000000000000000000000000111111110000000000000000000100000000000000000000000011110000000000000000000000000000000011110000000000001111000000010000000000000000000000000000000000000000000011110000000000010000111100000001000000000000000000000000000111110000000000000001000000000000111000000000000000000000000000000000000000010000000100000000000000000000000000001111000011111111000000000000000000000000000000000000111100000000000000000000000011100000000011111111000000010000",
		"00000001000000000000000000000000000000010000000000000000111100000001000000000000111100000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000011110001000000100000000000000001000000000000000000000000000100000000000000000001000011110000000000000000000000010001000000000000000000000001000100000000000000000000000000000000000000000000000000001111000000000000000100000000111100000000000000000001000011110000000000000000000000000000",
		"00010001000000000001000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000111100000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000011110001000000010000000000000000000000000000000000000000000000000001111100000001000000000000000000000000000000010000000000000000000100000010000011110000000000000000000000000000000100000000000000000000000000001111000000000000000000000000000011110000000000001111000000001111000000000000",
		"00010000000000000000000000000010000011110000000011110000000000000000000000000000000000010000000000000000000111110000000000000000000000000000000000000000000000001111000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000100000001000011111111000000000000000000000000000011110000000000000000000000001111000000000000000100000000000000000000111100001111000000000000000011110000",
		"00000000111100000001000000000001000011110001000000000001000011110000000000000000000000000000000000000000000000001111000000010000000100010000111100000001000000000000000000000001000000001111000000000000111000011111000000000000000000000000111100010000000000001111111100000000000000000000000000000000000000000000000000010000000000000000111100000000000000000000000000000000111100001110000000000000000000001111000000000000111100000000000000000000111100000000000000000000000000000000000000000000000000000000000011100001",
		"00000000000000000000000000001111000000000001000011110000000011110000000000000000000000011111000100000000000000000000000000001111000000000000111100000000111100000000000000000000000000000000111100000000111100000000000000000000000000000000000000010000000000001111000000000001000000000000000000000000000000000000000000000000000011100000111100000000000000000001000000000000000000000000000000000000000000000000000000000000000000001111000000000000111111110001000000000000000000001111000000000000000000000000000000000000",
		"00000000000000000000000000001111000000010000000000000000111100000000000000000000000100010000000000010000000000011111000000001111111100000000000000000000111100000001111111110000111100000000000000000000111100000000000000000000000000000001000000000000000000000000000100000001000000001111000000000000000000000000000111111111000011111111111000000000111100000000000000000000000000010000000000000000111100010000000000000000000000101111000000001111111111110001000000000000000011111111000100000000000000000000000000000000",
		"00010000000100001111111100011111000000001111000000001101000000000001000000000000000000000001000000010000000000001111000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000100000000000000000000011110000000000001111000000000000111111111110000000000000000011110000000011110000000000001111111100000000000000000000111100001111000100101111000100010001000000011111000000000000000000011111000000000000000011110001000000000000000011110000000000010000000000000001000000000000",
		"00000000111100011111000000001110000000001111000000011101000011110000000000001111001000000000000000100000000000011111000000011111000000000000000000000000000000000001000000010001000000000001000011110000000000100000000000010000000000000000000011110000000000001111000000000000000011111110000000000000111111110000000000000000000000001110000000001110111100000000111000001111000100010001000000000000000000001111000000010000000000000000111100000000111100000001000000000000000011110000000100000001000100000001111100001111",
		"00000000000000000000000000000000000000001111000100001111000000000000000000000000001011100000000000000000000000010000000100001111000000000000000000000000000000011111000000010010000000000001000100001111000100001111000000000000000100000001111011101111000000000000111100000001000000001111000100000001000000000000111100000000111100001111000000000000000011111111111100000000000100000001111100000000000000001111000000000000000000100000000000000000000000001110111100010000000000000000000000000010001000000000001000000000",
		"11111111000000000001111100001111000011111111000000000000111000000001000000010001000100000000111111110000111100000000000000000000000100011111111100001111000000011111000000010001111100000001000000010000000100101111000000000001000000000001111111110000000100000000000000000000111100011110001000000000000100000000000000010000111100000000000100001111111100010000000000010000000000010001111100010001111100000000111100000000000000010000000011111110000000001111000000001110111111110000111100000010000100000000001000001111",
		"00000000000100000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
		"00000000001000011111000000011111000000001111000100001111000000000000000111110000000011110000000100001111000011110000000011110000000000010001111000000000000100000001000000000000000000010000000011111111000000100000000000000001000000001111000000001110000111100001000100000001000100001111000000001110111100000000000111110001000000100001000000000000000000000000111100100000000000000000111100000000000000000001000100000000111111110001000100000001000000000001000000000001000100010000000000000000000100010000000000001111",
		"00001111000000000000000000001111111100000001000000001110000000000000000000000000000100000000000000000000000000000000111100001111000000001111000000000000000000000000000100010000000000000000000000001111000100010000000000000000000000010000000000000000000011111111000000010000000000000000001011101110111100000000111100010000000000010000000100001110000000001101111100000000000000000000000100011111000000000000000000000000000000000000000000000000000000000000000000010000000000000001000100000001000100001111000000010000",
		"00000001111100000001000000000000000000010000000100000000000000000001000000000000000100000000111100001111000011111110000000000000111000010000000100000000000000000001000000000000000000000000000100001111000000010000000011110000000000000000000000000000000011100000111100000000000000000000000111110000000000000001000000001111000000000001000011110000000000001111000000000001000000000000000111111111000000000000000000000000000000000000110100000000000000001111000000000000000100000001000011110000000000000001000000000000",
		"00000000000000000000111100000000000000000000000000000000111100000001000000000000000000000000111000010000111100000000000000000000000000000000000000000001000000010001111000010000000011111111000100000001111100100000000011110000111100000001000000000001000100000000000000000000000000000000000100001111111100000000000000001111111111110000000000001111000000000000000000000000000000010000000000001110000000000000000000000000000000000000110000000000111111110001111100000001000000000000000000000000000000000000000000010000",
		"00000000000000000000000000000000000011110000000000000000000011110001000000000000000000001111111000000000000000000000111100000000000000000000000000000000000000010001000000000000000011110000000000000000000000010000000000000000000000000001111100000000000111111111000000000000000000000000000000000000111111110000000000001111111100000000000000000000000000000000000000000000000000100000000000011110000000000000000000010000000000010000110100010000111011010001111100010000000000000000000000000000000000000001000000000000",
		"00000001000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000111100010000000000000000000100000000000000010000000000000000000000000000000000000000000000011111000000000000000000000010000000000000000000001111000000000000000000000000000000000000000011100000000000000000000011100000000000010000000100000000111100000000000000010000000000001110000000000000000000000000000000000000110000000000000011100000111000010000000100000000000000000000000100000000000011110000",
		"00000000000000000000000100010000000000000000000000010000000111110000000011110000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000001000000001111000100000000111100000000000011110000000000000001000000010000000000000000000000000000000100000000000011110000111111100000000000000000000011110000000000000000000000000001000000000001000000011110000000001111000000000000000000000000000000000000110000000001111111100000111100010000000100000000000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000101111000011111111000000001111000100000000000100000000000000000000000000000000000000000001000000000000000000000000000011110000000000000000000100000000111000000000000000000000000000000000000000001111000000000000000000000000000100000000000000000000111111110000000000000001000011111111000000000000000000000000000000000001000000001101000000011111000000000000000000000000000000010000110000000000000011100000111100000000000000000000000000000000000000000000000100010000",
		"11110000111111110000000000000000000000000000000000100000000000001111111111111111000100000000000100000000000111100000000000000000000000000001000000001111000000000000000011110000000000000000000100000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000100001000000000000000000000000000000001111000000000000000000001111000000000000000000000000110100010000000011110000000000000001000000000000000011110000000000001111000100100000",
		"00000000111000000000000000000000000000000000000000000000000000000000000000000000000100001110000000000000000111100000000000000000000000000001000000001110000000001111000011110000000000000000000000001111000000000000111100000000000000000000000100000000111100000000000000000000000000000000000000000000000000010000000000000000000011110000000000000001000000000000000000000000000000000000000100000001000000010000000000000001000000001111111100010000000011111111111100000000000000000000000000000000000000011111000000000000",
		"00001111110100000000000000000000000000000000000000000000000000000000000000000000000000001101111100000000000000000000000000000000000000010000000000001110000011100000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000100000000000000000000000000010000000000000000000000000000000000000001000000000000000000010000000000000000000000000000111100010000000000000000111100000000000000000000000000001111000000010000000000010000",
		"00010000111100000000000000011111000000000001000011110000000000000000000000000001000000001101000000000000000000000000000100000000000000001111000000000000000011110000000000001111000000000000000000001111000000000000000000000000000011110000000000000000000000000000000000010000000000000000000000000000000000011111000000000000111100100000000011110000000100000000000000010000000011110000000000000000000000000001000000000001000000000000000000000000000000001111111100001111000000010000111100000000000100100000000000000000",
		"00010000000000000000000000001111000000000001111000000000000000000000000000000001000000000000000011110000000000000001000100000000000000000000000000000001000011111111000100000000000000010000000000011111000000000000000000000000000011100000000000001111000000000000111100000000000000000000000011110000000000001111000000000000000000010000000011010000000100000000000000000000000111111111111100000001000000000000000000000000000000000001000000000001000000000000000000000000000000010001111100000001000100010000000000000000",
		"00000000000000000000000100000000000000000000111000000000000000000000111100000001000000000000000000000000000000000000000000000000000100000000000000000000000011110000000000000000000100010000000000000000000000000000000000000000000011110000000000100000000000000000000000000000000000000000000011110000000000000000000000000000111100000000000011100000001000000000000000010001000111111111000000000000000100001111000000000000000100000000000000000000000000000000000000000000000000000000111100000000000000000000000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000001000011110001000000000000000011110000000000000000000000000000000000000000000000000000000011111111000000000000000000010000000000010000000000000000000000000000000011110000000000100000000000000010000000000000000000000000000011110001000000000001000000000000111100000000000000000000000000000000000100000001000011111111000000000000000100001111000000001111000011110000000000000000000100000000000000000000000000000000111111110000000000001111000000010001",
		"00000001000000000000000000000000000000000000000000000000000000000001000000000000111100010000000000000000000000000000111100000000000000010000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000011110000000000010000111100000000000000000000000000000000000100000000111100000001000000000000000000000000000000000001000000000000000000000001000111110000000100000000000100001111000000000000000000000000000000000000000000000000000000000000000011110000000000000000000011110000111100010000",
		"00000000000000000000000000000001000000000000000000000000000000000000111100000000000000001111000000000000000011110000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000111100000001000000000000000000000001000000001111000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000001000000000000000000000000000011110001000000000000111100000001000000001111000000000000000011100000000000000000000000000000111100000000111000011111000000000001000000001111000000010000000000000000000000000000000011100000000000000000000000001111000000000000000011110000000011110000111100000000000000001110000000000000000000010000000000001111000000000001000011111111000000000001000000001111000000000000000000000000000000001111111100000000000000010001000000000000111100000000000000000000000000000000",
		"00000000000000000000111111110000000011110000000000000001000000000000111100000000000000000000000000010000000000001111111100000000000000000001111100000000111100010000000000000000111100001111000000010000000000000000000000000000111100000000111100010000000000001110111100000000000000000000000000000000000000000000000000001111000011110000111100000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001",
		"00000000000000010000000000001111000000000000000000001111000000000000000000000000000000001111000000000000000000001111000000010000111100000001111100000000111100000000000011100000111100000000111100000000111000000000000000000000000000000001000000000000000000000000000000000000000000000001000000010000000000000000000100000000000011100000111100001111000000010000000000000000000000000000000000000001000000000000000000000000000000001111000100000000000000000001000000000000000100000000000000000000000000001111000000000000",
		"00000000000000010000000000000000111100010000000000001110000000000000111100000000000000000000000000000000000000001111000000000000111100000000000000000000111100000001000011110000000000010000000000000000111000000000000000000000000011110001000011110000000000000000000100000000111100000000000000000000000000000000000111111111000000000000111000000000000000000000000000000000000100000000000000010001000000010000111100000001000000001111000000000000000011110001000000000000000000000000000100000000000011110000000000001111",
		"00010000000000011111111100011111000000001111000000001110000000000001111100010000000000000001000000000000000100001110000000000000111000000000000000000000111100000001111100000000000000000000000000000000000000010001000000000000000011110001000011100000000000000000000100000000000000000000000000001111111100000000001011111111000000001111000000001111000000000000000000000000001000000000000000010000000000010000000000000000000000000000000000000000000011110001000000000000000000000000000000010000000011110010000000000000",
		"00000000000000010000111100001110000000001101000000011111000000000000000000011111000100000000111100001111000000000000000000000000111100000000000000000000000000010000000000010010000000000000000100000000000100010000000000011111000000010001000011110000000000000000000011111111111100001111000000000000000100000000000100000000000000011111000011111110111111110000111000010000000100010000111100000000000000000000000000010000000100000000000000000000000000000000000011110000000000000000000100010001000100000001000000000000",
		"00001111000000000000000011110000000000011110000000001111111000001111111111110000001100000000000000000000111100000010000000001111111100000000000000000000000000011111000000010010000000000001000100010000000100001111000000001111001000000010111111100000111100001111000011111111000000000000000100000001000000000000000000000000111100001111000111110001000000000000000000000000000100010000111100000000000000000000000000100000000100010000000000100000111100000000000000010000111100010001001011110000001000000000001000000000",
		"00000000000000010000000000010000000000000000000000000000000000000010000000000001000000000000111100000000000000000000000000000000111000011111111000001111000000000000000000000000000000001111000000000001000100010000111100010001000100010001111111110000000011101111000000000010000000001111000100001111000000011111000000000000111000000000000000000000000000101110000000000001001000000000000000001111000011110000111111100000000100000000000000000000000000001111000100001111000000000001000011110001000000001111000000000000",
		"00000000000000000000000000000000000011110000111100000000000000000000000000000000000100000000000000000000000000000000111100000000000000001111111100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000011110000000000000001000000000000000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000011110000000000000001000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000010000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000",
		"00000000000100000000000000011111000000001111111100000000000000000000000111110000000000000000000000000000000011110000000000000001000000000000111100000000000000000001000000000000000000000000000000000000000000010000000000010001000000000000000000000000000100000000000100000001000000000000000000001110111100000000000000000001000000100001000000000000000000001111000100001111000100000000111100000000000000000001111100000000000000000001000000000000000000000001000000000001000000010000111100000000000000000000000000001111",
		"00001111111100010000000000001111000000000000000000001111111100000000000100000000000000000001111100001111000000000000000011110000111000000000000000000000000100000000000100010000000000010001000011111111000100010001000000010000000000010000000000000000000011111111111100000000000000000000000011111111111100010000000000010000000000010000000100001110111100001110111100000000000100000000000000001111000000000000000000010001000000000000000000000000000000000001000100010000000000000010000000000001000100000000000000001111",
		"11110001111011110000111100001111000000010000000000000000111100000000000000000000000000000001111100000000000000001111000000001111111100000000000000000000000100010001000000100000111100001111000000000000000100000000000011110000000000000000000000000001000011111111000011110000000000010000000000000000000000000010111100001111000000000001000000001111000000001111000000000000000000000000111100001110111100000000000100000000000000000000110111110000000000000000000000010000000000000010000000000000000000000000000000000000",
		"00000000000000001111111100011111000000000000000000000000111100000000000011110000000000000000111000000000111000010000000000001111111100000000000000000001000000100001111100100000000000001111000000000000111100010000000111100000111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111111111111000000000000000000000000000000000000000000010000000000001111000011110000000000000000000000000001111000000001111011100001000000100001000000000000000000001111000000000001000000010000",
		"00000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000111100000000111100000000000000000000000000010000111100000000000000010000000000110000000000000000000100000000111100000000000011100000000000000001111000000000000100000000000000010000000000000000000000000000000000000000000000010000111111110000000000000000000000000001111100000000000000011111000000000000000011111111000000000000000100000000111100000001111111110000111100100001000000000000000000000000000000000001000000000000",
		"00000001000011110000000000010000000000000000000000010000000000000001000011110000000000000000000000000000000000010000000000010000000000010000000000000000000000000000111100010001000000001111000000000000000000000000000011100000000000000010111100000000000100000000000000000000000100000000000000000000000011110000000000000001000011111111000000000000000000000000111100000000000000010000111100011111000100000000000000000000001000000000111100000000000011100000111000110001000000000000000000000000000000000000000100000000",
		"00000000000000000000000000000001111100000001000000000000000000001111000000001111000011110000000000000000000000010000000000000000000000000000000000001111000000010000000000010000000000000000000100000000111011111111000011110000000000000010000000010000000100000000000100000000000100000001000000000000000011010000111100000001000000001111000000000000000100000000000000000001000000001110111100000000000100010000000100000000000000000000111100000000000011110000111100100000000100000000000000000000000000000000000000000000",
		"11111111111100000000000000010000000000000000000000011111000100001111000011101111000011111111000100000000000100000000000000000000000000000001000000001111000000010000000000000000000000000000000000000000111000001111000000000000000000000001000000000000000000000000000100000000000000000000000000000000000011110000000000000001000000000000000000000000000100000000000000000000000000001111111100000000000000000000000000000000000100000000111100000000000011100000111100110000000000000000000000000000000000011111001000000000",
		"11110000111000000000000100000000000000000000000000011111000000000000000000000000000011111111000100000000000011100000000000000010000000000000000000001111000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000011110000111100000000000000000000000000010000000100000000000100000000000000000000000000000000000000000000000000000000000100001111000000000000000011110000111100100000000000001111000000000000000000001111000100010000",
		"00000000110100000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000011100000000000000010000000001111000000001111000000000000111100000000000000000000000000001111000100000000000011110000000000011111000011100000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000001000011110000000100000000000000000010000000000000000000010000000000000000000100001111000000000000000011111111111000010000000000000000000100000000000000011111000100000000",
		"00010000111100000000000000000000000000000000000011110000000000000000000000000001000100001101000000000000000000000000000000000001000000101111000000001111000000000000000011110000000000000000000000001111000100000000000000000000000100010000000000000000000000000000000000000000000000000000000000000001000000011111000000000000000000000000000000000000000011110000000000000000000000000001000000000000000100000001111100000000000000010000000000100000000000001111111100000000000000000000000100000000000000101111000000000000",
		"00010000000000000000000100001111000000000000111111110000000100000000000000000010000000001111000000000000000000000000000100000000000000001111000000000001000000001111000100000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011110001000000001110111100000000000000010000000011100000000011110000000000000000000011110000000000010000000000010000000000000000000000000000000000000000000000001111000000000000000000010000111100000000000000100000111100000000",
		"00000000000000000000000100000000000011110000111000000000000000000000000100000001000000000000000011110000000000000000000100000000000100000000000000000000111100000000000100000000000000010000000000001111000000001111000000000000000000000000000000001111000000000000000000010000000000000000000011110000000000000000111100000000000000010000000011010000000000000000000000010000000100001111000000000000000000010000000000000000000000000000000000000000000011110000111100000000000000010000000000000001000100010000000000000000",
		"00000000000000000000000000000000111100000000111100000000000000000000000000000001000000000000000011110000000000000000000011110000000000000000000000000000000000000000000000000000000000010000000100000000111100000000000000000001000011110000000000011111000000000000000000000000000000000000000111110000000011110000111100000000111100000000000011110000000100010000000000000000000100001111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001",
		"00001111000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000011110000000000000000000000001111000000001111000000000000000000000000000000000000000000000000000000000000000011110000000100010000000000000001000000010000000000010001000100000000000000000001000011110000000000000000000000000000000100000000000000000001000000000000000000000000000000001111000000000000000100001111000000000000000100001111000000010000000011110000000000010000000100001111000000000001",
		"00000000000000000000000000000001000000000000000000000000000000010000111100000000000000010000000000000000000011110000000000001111000000000000000000000000000000010000000000000001000000000000000000010001000000000000000000000000000111110000000000000000000000000000000100000000000000000000000000000000000000000000000000001110000000000000000000000000000100000000000000000000000100000000000000000000000000001111000000000000000000000000000000000000000000001111000000000000000011110000000000010000000000000000000000010000",
		"00000000000000000000000000000001000000000000000000000000000000000000111100000001000000001111000000010000000011110000000000010000000000000001000000001111111100000000000000000000000000000000000000000000111100000000000000000000000011100000000000000000000100000000000100000000000000000000000011110000111100000000000100001101000000000000000000010000000000001111111100000001000000000000000000000000000000001111000000000000000000000000000000001111000000001111000000000001000000000000000000000000000000000000111100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000010000111100010000111100000000000000010000000000000000111100000000000000000000111100000000000000000001000011110000000000000000000000001101000100000000000011100000000000000000111100000000000000001110000000001111111100000000000000011111111100000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000",
		"00000000000000000000111100000000000000000000000000000000000000000000111100010000000000001111000000000000000000000000111100001111111100000001111100000000000000100000000000010000111100000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000001111000000000000000100001111000011110000111000000000000000011111111100000000000000000000000000010000000000000000000000011111000000001111000000001111000000000000000000000000000000000001000000000000000011110000000000000000",
		"00000000000000010000000000001110000000000000000000001101000011110000000000000000000000000000111100000000000000000000000000010000111100010000000000001110000000010000000011110000111100000000000000000000111100001111000000000000000000000001000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000111100001111000000010000000000010000000000000000000000000000111100000000000000010000000100001111000011110000111100000000000000000000000000000000000000000000000011111111000000010000",
		"00000000000000000000000000001111000000000000000000001110000000000001111100000001000000000000111100000000000000000000000000000000000000000001000000000000000000000000000011110000000000000000000000000000000000000000000000010000000000000001111111110000000000000000000100001111000000001111000000000000111100000000000100001111000000000000000000000000000000000000000000000000000000010000000000010000111100000000000000000000000000001111000100000000000000000001000000000000000000000000000000000000000000001111000000000000",
		"00000000000000000000111100001111000000001110000000001110111100000001000000000000000000000000111100000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000111110000000000010000000000000000000011110001000011100000000000000000001000000000000000000000000000001111111111100000000111110000001000010000000000000000000000000000000000000000001000100000000000010000111100000000000000010001000011110000000000000001000000000000000000000000000000010000000100000000000000000000000000000000",
		"00000000111100001111111100011111000000001101000000011111000011110000000000000000000000000000111100000000000000000001000000000000111100000000111100000001000000000000000000000001000000000001000100001111000100000001000000100000000000010001000011100000000000000000000000000000111100000000000111110000000011110000001011010000000000010000000011110000111111110000000000000000000000100000111100010000111100000000000000010001000011110000000000010000111100000001000011110001000000000000000000000001000000010000000000000001",
		"00011111000000000000000011111111000100011110000100000000111000011110000011100001001000000000111100000000000000010010111100001111111000001111111100001110000000010000000000010010111100010001000100011111001000001110000000000000001100010001111011101111000000000000000000000000111100001110001100000010000011111111000011110000111100000000000111110001000000000000000000100000000100110000000000001111000011110000111100010000000000010000000000011111111000001111000100001111111000000000001000001111010000001111001011110000",
		"11111111000000000001000000001110000000000000000000011111000000000010000000000001000000000000111011110000111100000000000000001111111100001111111000000000000000011111111100010001000000000000000100000000000100110000111100010000000000000010111111110000000011110000000000000000000000001110000000000000000000000000111100000000111000000000000100000000111100000000000000010000001000010000111100000000000011110000111011110000000100001111000000001111000000001111000000011110111111110000000000000010000100001111000100001111",
		"00000000000011110000111100000000000000000000000000000000000000000001000000010000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000111100000000000000010000000000000000000100000000000000000000000000000000000000010000000000000010000000000001000000000000000000001111111111110000000000000000000000000000000000010000000011110000000000000000000000010000000000000000000000000000000000000000000000001111000000010001000000000000001000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000100000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000001000000010000000011110000000000001111000000010001000000000001000000000001000000000000000000000000000100000001111100000000000000000000000000000000000000010000111100010000000000000000000000010000111100000001000000000001000000000000000100001111001000000010000000000000000000000000111000000000000011110000000000010000000000010000000000011111000000000000001000000000111100010000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000011110000000000001111000000001111",
		"00001111111100010000111100001110000000001111000000001111111100010000000000010001000011110000111100000000111100000000000011110000111100000000111000000000000000000001000000000000111100000001000011110000000000000000000000001111000000000000000000000000000011111111111111110000000000001110000000000000000000101111000100100000000000010001000000001110111100001111000000000000000000000000000000010000111100000000000000010000000000000000000011110000000000000000000100000000000000010001000000000001000000010000000011110000",
		"00000000111000000000111100000000000000010000000000000000111100000000000011110000000000000001000000001111000000000000000100001110000000010000000000000000000000000000000000100000000000000000000011110000000000000000111111110001000000000000000000000000000000000000000011110000000000001111000011110000111100000000111100100000000000000000000000000000000000001111000000000000000100000000111000000000111100000000000000000001000111110000000011110000111100000000000000010000000000000001000000000000000100000000000000010000",
		"11110001000000000000111100001111000000000000000000000000000000000001000000000000000000000000000000001111111000010000111100001110111100000000000000000000000000010000111100100000000000000000000000000000000000000000000011010000111111110000000000000000000000000000000100000000000000001111000100001101000000000000000000001110000011111111000000000000000000000000111100000000000000010000000000001111111100000000000000000000000000000000000011110000111100000000000000010001000000000000000100000000000000000001000000010000",
		"00000000111100000000000000011111000011110000000000100000000000000001000000000000000000001111111100000000111100000000000000001110000000000000000000000000000000010000000001000000000000000000000000000000111000000000000011010000111100000000111100010000000000000000000000000000000000000000000000001110000011110000000000001111000011111111000000000000000000000000111100000000000000011111000000000000000011111111000000000000000100000000000000000000111111110000000000100001000011110000000000000000000000000001000000010000",
		"11110001111100000000000000000000000000000000000000100000000000000010111100000000111100001111000000000000000000000000000000001111000000000001000000000000000000010000000001000001000100000000000000000000111100000000000011100000000000000000111100000000000000000000000000000000000000000001000000000000000011110000000000000000000000000000000000000000000000000001111100000000000000011111111100000000000000001111000100010000001000001111000000000000000011100000111100110001000000000000000000000000000000000000000000000000",
		"11110000000011110000000000000001000000000001000000000000000000000000000011101111000000000000000000000000000000000000000000000000000000010000000000001111000000010000000000110001000011110000000000000000111000001111000011100000000000000001000000010000000011110000000000000000000100000001000011110000000011100000000000000000000000000000000100000000000000000000000000000001000000011111000000000000000100000000000100000000000100000000000100000000000011110000000000100001000000000000000000000000000000000000000100000000",
		"11100000111111110000000000000000111100000001000000010000000000001111111100001111000111111110000100000000000000000000000100000000000000000000000000001111000000010000000000110001000100000000000000000000111011110000000011100000000000000000000000000000000100000000000100000000000000000001000000000000000111010000111100000000000000000000000100000000000000000000000000000000000100000000000000000001000100010000001000000000000100000000000000000000000011110000111100110000000100000000000100000000000000000000001000001111",
		"11100000110111111111000100000000000000000000000000000000000000000000000000000000000100001110000000000000000000001111000000000001000000000000000000001111000000100000111100010001000000000000000100000000000000000000000011110000000000000000000011100000000100000000000000000000000000000001000000000001000011010001111000000000000000000000000100000001000011110000000100000000000000000010000000000000000000000000000000000000000000000000000000000001000011111111111100100000000000000000001000000000000000000000001000000000",
		"00000000111000000000000100000000000000000000000011110000000000000000000000000000000100001110000000000000000011111111000000000001000000000000000100000000000000010000111100010001000000000000001000000000000100000000000011110000000000000000000011110000000000000000000100000000000011110000000000000000000011110000111000000000000000010000000100000000000000000000000000000000000000000010000000000000000100010000000000000000000000000000000000000000111111110000111100101111000000001111000100000000000000010000000000000000",
		"00010000000000000000000100000000000000000000000011110000000100000000000000000001000000001110000000000000000000000000000100000001000000001111000000000001000000000000000000010001000000010000000000000000000111110000000011110000000100000000000000000001000100000000000000001111000000000000000011110001000000000000111100000000000000010000000011110000000011010000000000000000000100000010111100000000000000000000111100010000000000000000000000000000111111110000111100101111000000001111000000000000000000011111000000000000",
		"00010000000000000000000100000000000000000000111111110000000000000000000100000000000000000000000011100000000000000000000100000001000000001111000000000000000000001110000000010000000000000000000000010000000000001111000011100000000000000000000100000000000000000000000000010000000000000000000000000000000000000000111000010000111100010000000011100000000011110000000000010000000100000000000000010000000000000000000000000000000000000000000000000000000000000000111100010000000000010000111100000000000100011111111000000000",
		"00000000000100000000000100000000000000000000111011110000000000000000000000000000000000000000000111100000000000000000000000000000000100000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000100000000000000000000000000000000111100000000111100000000000011110000000000010000000000010000000000000000000000000000000000000000000100000000000011110001000000000000000011110000000000000000000000000000000000000000000100000000000000000000",
		"00000000000100000000000100000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000011110000000000000000000000000000000000000000000011100000000000000000000000000000111100010000",
		"00000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000001111000000010000000000000000000100000000000000010000000000000000000000001111000011111111000000010000000011110000000000000000000000000000000100000000000000000000000000001111000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000011111000000000000000000000000",
		"00000000000000000000000000000000111100000000000100000001111100010001111100000000000000000000000000010000000011110000111100010000000000000001000000000000000000100000000100000000000000000000000000000000000011110000000100000000000011110000111100010000000000001111000000000000000000000001000000000000000000000000000000001110000000000000111100010000000000001111000000000000000000001111000000000000000000010000000000010000000000000000000011110000000000000000000000000000000000000001000000000000000000000000000000000000",
		"00001111000000000000000000000000000000000000000000000001000000000000111100000000111100000000000000000000000000000000111100100000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000001000011110000111100000000000100001110000100010000000000000000000100001111111100000000000000001111000000000000111100010000000000100000000000000000000000000000000000000000000100010000000000000000000100000000000011110000000000001111000000000000000000000000000000000000000000010000000000000000",
		"00000000000000001111000000000000000000000000000000010000000000000000111100000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000111100000000000100001101000000000000000011110000000000000000111100001111000100000000000000010000111100000000000000000000000000000000000000010000000000000001000100001111000000011111000000000000000011110000111100000000000000000000000000000000000000000000000000011111000000000000",
		"00000000000000001111000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000000000000000011110000000100000000000000000000111111110000000000001111000000010000000011110000000000001111000000000000000000000000000000000000111100000000000000010000111100001111000000010000000000000000000000010000000000011111000011110000000000000000111100000000000000001111000000000000000000000000000000001111000000000000",
		"00010000000000010000000000001111000000000000000000001101000000000000000000000000000000000000111111110000000011110000000000000000000000010000000000001111000000011111000000000000000000000000000000001111000000000000000000000000000000000001111100000000000000000000000100010001000011111111000000000000000000000000000011110000000100000000000000000000000000010000000000001111000000010000000000000000000000010000000000011111000011110000000000001111111100000000000000000000000000000000000000000000000100001110000000000000",
		"00010000000000001111000000001111000000000000000000011110000000000001000000000000000000000000000000000001000100000000000000000000000000010000000000000000000000000000000000000000000000000000000011110000000000000000000000000000111100000000111111110000000000000000001000011111000000000000000000001111000000000000000111110000000100100000000000001111000000000000000000001111000100000000000000010000111100000000000000010000000000000000000000001111000000000000111100000000000000000000000000000000000000000000000011100000",
		"00000000000000000000000000000000000000000000000000010000000000000000111100000000000000000000000000000001000000000000000000000000000100000001000000000001000000000000000000000001000000010000000011111111111100000000000000000000000000000010000000000000000000000000000100000000000011111111111100000000000011110000000011100001000100011111000100000000000000000000111100000000000100000001000000000000000000000000000000000000000000000000111100010000000000000000000000000001000000000001000000000000000000010001000000000000",
		"00010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000010000000100000000111100000010000000000000000000000001000000000000111100000000000011110001000000000000111100000001111100000000000000000000000100000000111111110000000000000000000011100000000011100010111100000000000000010000000000000000111100000000000000000001111100000000000000000000000000000000000000000000000000000000000000011111000000000000111100000000000000010001000000100001000000000000",
		"00010000001011110000000000000000000000000000000000000000000011110000000100000001000100001111111100000000000000010000000000101110000000010000111100001111111100011111000011110000111100001110000100010000000100001111111000010001000000010000000011110000001000010000000100010000000000010000000100000001000011100001000000000010111100000000000000000000111100010000000000101111000111110001000000000000000011110000000011100000000000010000001000001111111000010000001000011110111011111110000000000000000000000000001100010000",
		"00000000000100000000000000010000000000000000000000000000001000000010000000010000111100000001111111110000000011111111000100000000001011110000000000000001111100011111111100000000111100001110000000000000111111110000000000010001111100000000111100000000000000000000000000000000000000000000000000000001000100010000111100000001111000000000000000000000000000000000000000000000000011110001000000000000000000001111000011100000000000000000000011111111000000101111000000011111000000001111111100100001000000000001000111110000",
		"11110001000100000001111100000000000000000000111100000000111100000001000100011111000111110000111000001110111111111111111100010000001011110001111100000000001000000000000000010001000111100000000111110001000111110001000000010000111000000000111100000001001000000000000000001111000000010001000000000001000000000000000000010000000000000000000000011111111111100001000011110000001000010000000011100001000011100000000011100001000000011111000000000000000000010000000000000001000111111111000000010010000000000001001000001111",
		"00000000000000000000000000000000000011100000000000000000000000000000000000000000000000000001000000000000000000001111000000000000000100000000000000000000000000000000000000000000111111110000000000000001111100000000000000000000000000000000000000000001000000000000111100001111111100010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000010000000000001111111100000000111100000000111100000000000000000000",
		"00000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000011100000000000010001000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000010000000000010000000011110000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000100000000000000010000000000000000000000000000000000000000000000000000000000000001000000001111000000001111000100000001000000000000000000000000000000000000000000000000111100000000000000000000111100000000000000000001000000000000000000000000000000001111000000000001000000000000000000000000111100000000000000000000000000010000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000001111000000000000000100000000000000000000000000000000000000000001000000000000111111111111",
		"00000000111000100001111100011111000000000000000000001110111000100000000000000011000000000000000000000000000000000000000011110000111100000000111000001111000000000001000000000000111100000000000000000000000000001111000000000000000100000000000000000000000011100000000000000000000000001110000011110000111000101111000100010000000000010000000000001111000000001110000000000000000100001111000000010000000000000000000000000000000100000001000111111111000000000000000011100000000000010000000011110000000000001111000000000000",
		"00000000000000010000111100000000000000000000000100010000111100000000000100000000000000000000111100001111111100000000000000000000111100000000000000001111000000000000000000010000000011110000000000001111000011111111000000000000000000000000000000000000000000000000000000000000000100001111000000000000111100001111000000000000000000011111000000001111000000001111000000000001000000010000000000000001000000000000000000000001000000000000000111101111000000000000000000000000000000000000000000000001000000000000000100010001",
		"00000001000000000000000000001111000000000000000000100000000000000001000000000000000000010000111111110000111100000000111100001110000000000000000000000000000000000000000100010001000000000000000000000000000000000000000011100000000011110000000000010000000000000000000000001111000000001110000000001110111100001111000000011111000000001111000000000000000000010000111100010001000000101111000000000000111100001111000000000000000111110000000011110000000000000000000000000000000000000000000100000000000000000001000000000001",
		"11110001000000010000000000000000000000000000000000010000000000010001000011110000000100101111000000000000000000000000000000001101000000000000000000000000000000000000000000100001000000000000000000000000111000000000000011100000000011110000111100010000000000000000000000000000000000001111000000001110000100001111000000001110111100000000000000000000000000000000111100000001000000101111000000000000111111111111000000100000000000010000000100000000000000000000000000000001000000000001000111111111000000000000000000000000",
		"00000000000000000000000000000000000000000000000000010000000000010000000011110000000100001110000000000000000000000000000000001101111100000000000000000000000000010001000000110000000000001111000000000000110100000000000011110000000000000000111100010000000100000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000101111000000000000000000001111000100010000000000001111000000000000111100000000000000000010000000000001000000000000000000000000000000000000",
		"00000000111100000000000000000000000000000000000000000000000000000000111100000000000100001111000000000000000000010000000000001100111100000000000100001111000000010000000000110000000011110000000100000000110100000000000011110000000011110000111100010000000100000000000000000000000100000000000000000000000011110000000000000001000000000000000000010000000000000001000000000001000000101111000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000100000000000000000000000000000000",
		"11110000111100000000000000000000111100000001000000000000000000000000000011110000000100001101000100000000000000010000000000011110000000000000000000000000000000010000000001010001000000001111000000000000111100000000000011100000000000000000000100000000000100000000000100000001000000000000000000000000000011110000000000000001111100000000000000000000000000000001000100000000000000100000000000000000000000000000000100000000000000000000000100000000000000000000000000010000000000000000000100010000000000000000001000000000",
		"00000000111011110000000000000000000000000001000000000000000000000000000000000000000100001101000000000000000000000000000000001111000000000000000000000000000000010000000001000001000000010000000100000001001000000000000111010000000100000000000011110000000100000000000011110000000000000001000000000010000011100000000000000001000000010000000100000000000011110001000100000000000000010010000000000000000000000000000000000000000100001111000000000000000000000000000000010000000000001111000100000000000000010000000100000000",
		"00000000111111110000000100000000111100000001000011110000000000000000000000010001000000001110000000000000000000000000000000000000000000000000000100000000000100010000000000110001000000001111000100000000001000000000000011010000000100000001000000000000000000000000000011111111000011110000111100000010000011100000111100100001000000000000000011110000000011110000000000000000000100010001000000000000000100000000000000000000000000000000000100000000000000000000000000010000000000000000000111110000000000000000000000000000",
		"00100000000000000000000000000000111100000000000011110000000100000000000100000001000000000000000000000000000100000000000000000000000000000000000100000001000000101111000000110001000000001111000000000000000100000000000011000000000000000000000000010000000000010000000000001111111100001111000000000001000011101111111100100001111000010000000011110000000011110000000000010000000000010001000000000000000100010000000000010000000000000001000100000001000011110000111100010000000000001111000100001111000100010000111000000000",
		"00100000000000000000000000000000000000000000111111110000000100000000000000000000000000010000000011100000000100000000000100001111000000001111000000000000000000011111000000010000111100001111000000000000000000001111000011000000000000000000000000000000000100000000000100010000000000000000000000000001000000000000000000000000111100000000000000000000000000000000000000010000000000010000000000010000000000000000000000010000000000000000000100000000000011110000111100000000000000000000000000000000000000000000111100000000",
		"00000000000100000000000000000001111100000000111000000000000100000000000000010001000000000000000011100000000000000000000000001111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011110000000000000000000100000000000000000000000000010000000100000000000000000000000000000000000000000000111100000000000000000000000000100000000000010000000000000000000100000000000000000000000100000000000000000000000000000001000011110000000000000000111100001111000000001111000100000000000000000001",
		"00000000000111110001000000010000000000000000111100000000000000010000000000000000000000000000000000000001000000000001000000001111000000000000000000000000000000010000000000010000000000000000000000100000000100000000111100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001110111100000000000000000000000000010000111100000000000000000000000000000000000000000000000000000001000011110000000000000000000000000000000000010000000011110000000000011111000000000000111100000000",
		"00000000000000000000000000010000000000000000000000000001000000010000000000000001000000000000000000010000000000000000000000001111000000000000000000001111000000010000000100000000000000000000000000010000000000000000111100010000000000001111111100000000000000001111000000000000000000000000000100000000000000000000000100001110000000000000000000010000000000000000111100010001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000",
		"00000000000000000000000000010000000000000000000100000010111100010001000000000000000000000000000000010000000000000000111100010000000000000000000100000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000111100000000000000001111000000001111000000000000000100000000000000000000000000001111000000000000000000000000000000010000000000010000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000111100000000",
		"00000000000000000000000000010000000000000000000000000000111100010000000000000000000000000001000000010000000000000000000000010000000000000000000000000000000100010000000000010000000000000000000000000001000000000000000100000000000000000000000000000000000100001110000100010000000000000000000000000000000000000000000000000000000000000000111100010000000000010000000000010000000000010000000000000001000000000000111100010000000000000000000011110000000000000000000000000000000000000000000000010000000000001111000000000000",
		"00000000111100000000000000000000000000000001000000010000000000000000000000000000000000000001000000000000000000000000111100010000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000100000000111100000000000000000000000000001110000000011111000000000000000000000000000000000000000000000000000000000000111100000000000000010000000000000000000000101111000000000000000000000000111100010000000100000000000011111111000000000000000000000000000000000001000000000000000000001111000000000000",
		"00000000000000011111000100001111000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000001000000001111000000000000000100000000000000000000000000001111000000001111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111100001111000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000010000",
		"00000000000000010000000000000000000000000000000000001110000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000001111000000000000000100000000000000010000000011111111000000000000000000000001111100000001000000000000000000000001000100010000000000001111000000000001000000000000000000000000000100000000000000010000000000011111000000001111000100010000000000000000000000000000000000010000000011110000000000001111000000000000000000000000000000000000000000000000000000001111000000000001",
		"00000001000000000000000000001111000000000000000000011110000000010000000011110000000011110000000000000000000000000000000000000000000000010001000000000000001000000000000100000000000000000000000000000000000000000000111100000000000000000001111000000000000000000000000000000000000000001111000000000000000000000001000000000001000100100001000100000000000000001110000000001111001000010000000000000000111100000001111100010000000000011110000000001110000000000000000000000001000000000000000000000001000000000000000000000000",
		"00000001000000000000111100000000000000001111000000101111000000010000000000000000000000000000000000000001000000000000000000000000000100010000000000000000001000000000000000010000000000010001000000000000000000000000000000000000000000000010111100001111000000001111000011110000000000001110000000000001000011100000000000000001000000101111000100011111000000001110111100001111000100010000111100000000111100000001000000010000000000011111000000001111000000001111000000000010000000000000000000010000000000100010000100000000",
		"00000000000000000000000000000000000000000000000000010000000000001111000000000000000000000000000000000000111100000000000000001110000100000000000000000000000000010000000100010001000000000000000000000000000011110000111100001111000000000001111100000000000000001111000000000000000000001110000100001110000011100000111111010001000000100000000000001111000000000000000000010000000100000000000000000000000011110000000000010000000000101111000000000000000000010000000000001110111111111111000100000000000000010001000100000000",
		"00001111000000000000111100100000000000001111000000000001000000000000000100000000000100001111111100000000000000100000000000010000000100000000111100000000000000011111000000000000111100001111000000000000000000000000000000000000111100000000000011110000001000010000000000000001000000000000000000000001000000000001000000000010000000100000000111100000111100010000000000101111000000000000000000010000000011110000000000000001000100010000000000000000111100000000000000001110111000001101000011110000000000010001000100000001",
		"00100001000100010000000100010000111100000001111100010000001011110010000000010000000000000010111111110000000011111111000100000000001000000000000000000001111100011111000011111111111011111110000000000001111011110001000000000000111100000000111100100001000000000000111100000000111100000001000000010000000000000010111000000001111100000000000000000000000000000000000000000000000011110001111100000001000000001110000011100010000000000001000111110000000000100000000000010000000011111111111100010001111100000010000100010000",
		"00001111000100000000000000000000000000000001000000000000000000000000000100000000000000000001000000001111000011110001000000000000000000000000111100000000000000000000000000000000000000000000000100000000000000000000111100010000000000010000000000000001000011110000000000000000000000010000000100000000000000000000000000000001000000010000000100000000000000000000000000000000000000000000000000000000111111110000000000000000000000010000000000000000000000001111000000001111000011110000000000000001000100000000000100010000",
		"00001111000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000111100001111000000000000000000000000000000010000000000000000000000000000000000000000000011110001000000010001000000000000000000000000000000000001000000000000000000000001000000000000111100010001000000000000000000010000000000000000000000000001000000000000000000000000000000000001000000000000000011110000000000000000000000000001000000000000000011110000",
		"00000000000000000000000000000000000000000000000000010000000111110000000000001111000000000001111100000000000100001111000000000000000000000000000011110000000000010000000000001111000011110000000011110001111100000000000000010000000000000000000000000000000000011111111100000000000000000000111100000000000000000000000000000000000000000001000000000000000000000000111111110000111111110000000000010000000000000000000011110000000000001111000000000000000000010000000000010000000000000000111100010000111100000001000000000000",
		"00000000000100000000000000000000000011110000000100000000000000000000000000000000000000000000000000000000000000000000111100000001000000010000000000000000000000000000000000000000111100000000000000000000111100000000111100010000000000010000000000000000000000000000000000000000000000000001000000000001000000000000000100000000000000000000000000001111000000000000111100010000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000100000000000011110000000000000000000000000000111111110000",
		"00000000000000100001111000001111000000000000000100000000111000000000000000100001000000001111000000010000000100000000000011110001111000000000111100001111000100000000000000000001000000000000000100001111111100010000000000000010000000000000000000001111000011111111000100000001000000001111000011111111111000010000000100000000000100011111000000000000000000001110000000000001000100001111111100000000001000001111000011110000000000000001001000001111000000000000000011110001000000000000000000000000000000000000111000000000",
		"00000000000000000000000000000000000000000000000100010000111000010001000000000000111100001111111100010000111100000001000011110000111100000000000000000000000000000000000000000001000000000000000011110000000000001111000000000000000000000000111100000000000000001111000100001111000100001111000000000000000000000000000000000000000000000000000000000000000000001111111100000001000000000000000000000001000011110000000000000000000000000000000111101111000000000000000000000000000000000000000000010000000000000000000000000001",
		"11110000111000000000000000000000000000000000000000010000111100000001000000000000000000000000111100000000111100000000000011111110111111110000000000000000000000000000000000000001000000000000000100000000000000000000000011110000000000000000000000000000000000001111000000000000000000000000000011111111000000001110000000000000000000000000000000000000000000000000000000000001000000010000000000000000000011110000000000000001000000000000000100001111000000000000000011110000000000000010000100000000111100000000000000000000",
		"00000000000000010000000000000000000000000000000000000000000000000001000000000000000000011111000000000000000000000000000000001101000011100000000000000000000000000000000000010000000000000000000000000000111000000000111111110000000000000000000000011111000011111111000000000000000000001110000000001101000000001111000011100000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000010000000000000000000100001111000000000000000000000000000000000001000111110000000000000000000011110000",
		"11110000000000000000000000010000000000000000000000000000000000000000000000000000000000001110111100000000000000000000000000001100000011110001000000000000000000000000000000100000000000000000000000000000111000000000000000000000000000000000111000001111000000000000000000000000000100001111000000001111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000111110000111100000000000011110010000000000000000000000000000000000000000000000000",
		"11110000000000000000000000000000000000000000000000000000000000010000000000000000000000001110111100000000000000000000000000001011111111110000000100000000000100000000000000010000000011110000001000000000101100000000000011110000000011110000111000010000000000001111000011110000000100001111000000001111000000000000000000000000000000000000000000011111000000000000000000000001111100100000000000000000111100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000100000000",
		"11110000111100000000000000010000000000010000000000010000111100010000000000000000000000001110000000000000000000000000000100001010000011100000000000000000001000000000000000010000000000001111000100000000111100000001000011110000000000000000000000000000000100010000000000000001000000001111000000000000000000001111000000000010000000010000000000001111000011110000000000000000000000100000000000000000000011110000000000000000000000000000000100000000000000000000000000000000111100000000000000000000000000011111001000000000",
		"00000000111100000000000000000000000000000001000000000000000000010000111100000000000000001111000000000000000000000000000000001001000011100000000000000000001000000000000000100001000000011111000100000000000100000001000111110000000011110001111111110000001000010000000000000000000000001110000000010000000000000000000100000000000000001111000011110000000011100001000100000000000000010001000000000000000000000000000000000000000000010000000000000000000000000000000000000000111100000000000100000000000000010000000111110000",
		"00010000000000000000000000000000111100000000000000000000000000000000000000000001000000011111000000000000000100010000000000001011111111100000000000000000000000010000000000100001000000011111000000000000000000000000000000000000000100000001000000000000000100000000000000000000000000001111000000000001000000000000000000000001111100001110000011110000000011110000000000000000000000010010000000000000000000001111000000000000000100000000000000000000000000000000000000000000000000000000000011111111000100000000111000000000",
		"00010000000100000000111100000000000000000000000100000001000000000000000000010000000000010000111100000001000100001111000000001101000011100000000000000001000100010000111100100000000000001111000000000000000000000000000011101111000000000000000000000000000000010000000000001111111100000000111000000000000000000000000100010001111100000000000011110000111111100000000000010000000000100000000000000000000000000000000000010000000000010000000100000000000000000000000000010000000000000000000000000000000000000000111000000001",
		"00010000000100000000000000000000000000001111111100000000000000000000000100000000000000010000111111010000000100000000000000001101000011100000000000000000000100001111111100010001000000001111000000000000000000001111000011100000000000000000000000000000000000000000000000000000000000000000111100000000000000010000000100000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000100100000000100000000000100010000000000000000000000000000000000001111000000000000000100000000000000000000",
		"00000000000100000000000000000001111111110000111100000000000000010000000000000001000000000001000011110000000100000001000000001111111111110000000000000000000000010000111100000000000000001111000000000000000000000000111100000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100001111111100000000000000011111000000100000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000100000000000000001111000000000000000100000000000000010000",
		"00000000000000000000000000000000000000000000111100000000000000010000000000000001000100000000000100010000000011110001000000000000000000000000000000000000000000010001000000010000000000001111000000010000000100000000111100010000000000000000111100000000000000001111000000000000000000000000000100000000000000010000000100001111000000000000000000000000000000100000000000010000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000010000000000000000000000000000111100010000000000000001000000000000000100100000000000000001000000000000000000000000000000000000000000000000000100010000000000010000000000010000000000010000000000010000000100000000111100000000000000000000000000000000000100000000001000000000000000000000000000001111000000000001000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00001111000000000000000000001111000100000001000100000000111100000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000100000000000000001111000000000000000000000000000000000000000000000000000000001111000000010000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000111100000000",
		"00000000000000000000000000000000000100000001000100000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000011111000000000000000000000001000000000000000000000000000000001111000000000000000000000000000000000001000000000000000000001111000000000000",
		"00000000000000000000000000000000000000000001000000011111000000000000000000000001000000000000000000000001000000000000000000000000000011110000000000000001000100000000000000001111000000000000000000000000000000000000000100000000111100000000000000000001000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000011111000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001110000000000000",
		"00000000000000001111000000000000000000000000000000101101000000010000000000000000000100000000000000010000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000011111111000000000000000000010000000000000001000000000000000000000000000000010000000100000000000000000000111100000000000000000000000000000000000000000000000000011111111111111111000000010000000011110000000000000001000000010000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
		"11110000000000000000000000000000000000000000000000001101000000100000111100000000000000000000000000000000000000000000000000000000000000000000111100000000000111110000000000000000000000000001000011111110000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000001111100000000000000000000000100010000000000000000000000001111000000000000000000000000000000000000000000000000000000010000000000001111000000000000000000000000000000000000000000000000000000010000000000000000000100010000",
		"00000000000011110000111100001111000000001111000000011110000000100000111100000000000000001111000000000000000000000000000000000001000000000001000000000000000100000000000100010000000000000000000000001111000000000000111100000000000011110001000000000000000000000000000000001111000000001111000000000001000011110000000000000000000100100000000000000000000000001110000000001111000000010000000000000000111100000001000000010000000000101110000000001111000000001111000000000001000000000000000000000000000000010000000100000000",
		"00000000000000000001000000001110000100000000111100011111000000100000000011100001000000000000000000000001111100000001000000000001000000000000000000000001000111110000000100000000000000000010000000010000111100000000111100001111000100000001000011110000000011110000000000000000000100001111000100000000000011110000000000000001000000110000001000000000000000000000000000000000000000100000111100000000111011110001000000100000000000111111000100001111000000001111000000000001000000000000000000000000000000010001000100000000",
		"00000001000000010000000000001111000000001111000000010000000000000000000000000000000000000000000000010000000000000000000000001111000100000000000000000001000000000000000000101111000100000000000000000000000000000001000000001111000011110000000000000000000000000000111100010000000111111111000000001111000000000000111100000000000000000001000000000000000000010000000000000000000000100000000011111111000011110001000100010000000000000000000011110000000000010000000000001110000000001111000011110000000000000010000000000001",
		"00001110000100001111000000100000000000001110000000010000001000001110000011110000000111110000111100000000000000010001000000000001000000010000111100000000000000001111000000001111000000000001000100001111000000010000111100000000111100000000000011110000000111110000000000010000000000000001000011110000111100000001111100000010111100100001000111100000111000100000000000111111000000000000000100011111111111110010000011110000000100000000000011110000000000000000000011111110111000001101000111110000000000010001000000000000",
		"00000000000100000001000000011111000100000000000000000000000000000000000000000001000111110010111111111111000000000000000000000000000000011111111000000000000000001111000000010000000000000000000100000000000100000000111100000000000000000001000011110000000111110000000000000000000000000000000000011111000000000001000000000000000000000001000100001111111100000000000000010000000100000000000000000001111111110001111111110001000000000000000000000000000000001111000000000000111111110000111100000001000100010000000000000000",
		"00000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001111000000000000000000010000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00001111000111110000111100000000000011110000000000000000000000000000000100000000000000000000000000001111000011110000111100010000000000000000000000000000000100000000000000000001000000000001000100000000000000000000111100000000000000010001000000000000000000001111000000000000000000000000000000010000000111111111000100000000000000010000000000010000111100010000111100100000000000000001000000000001000000000000000000000000000000010000000100000000111100001111000100010000000000000000000100010000000100000000000011110000",
		"00000000000100010001111000001110000000001111001000011111111000010000000100000010000000001111000000001110000111110000000000000001111000000000111000001111001000000000000011110001111100000000000100001111111100010000111000000001000000000000000000010000000011100000000100000001000000000000000000000000000000000000000000000000000000010000000000000000000000001110000000010001000100000000111100000001000100000000111111110001000100000000001000001110111100001111000111110000000011110000000000000000000000000000000000000000",
		"11100000000011110000111100000000000100000000000000000000101100000001000100000000000000001111111100010000000000000000000000000000000011110000111100001111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100010000111100000001000000000000000011110000000000010000000000000000000011111111000000000000000000000000111100000000000011110001000000000000000000011111000111101110000000000000000000000010000000000000000000010000000000000001000100000001",
		"11110000111100000000000000000000000100001111000000000000111000000001000011110000000000001111000000010000000000000001000000001111111111010000000000000000000000001111000000000000000011110001000000010000111100000000000000000000000011110000000000010000000100000000000000000000000100010000000000000000000000000000000011110000000100000001000000000000000000000000000000000001000000000000000000000000000011110000000000000000000000000000000000000000000000010000000011110000000000000000000000000000111111110001000000000000",
		"11110000000000010000000000010000000000001111000000000000000000000000000100000000000000000000000000000000000000000000000000001110000011100001000000000000000000000000000000001111000000000001000000000000111100000000000000000000000000000000111100001111000011110000000000000000000100000000000000000000000000000000111111100000000000000001000000001111000000010000000000000001000000000001111100000000000011110001000000000000000000000000000100000000000000000000000111110000000000010000000000000000111100000001000011110000",
		"00000000000000000000000000100000000000000000111100000000000000000000000011110000000000001111000011110000000000000001000000001110000011100001000000000000000000000000000000000000000000000000000000001111110000000000111100000000000000000000111000000000000100000000000000000000000000001111000000001110000000010000000011110000000000000000000000000000000000000000000000000000000100000000111100000000111100000000000000000001000000000000000000001110000000000000000000000000000000010000000000000000000000010000000111111111",
		"11110000000000010000000000000000000100000000000000000000111100000000000000001111000100001110000000000000111100000000000000001101111111100000000000000000000100010000000000000000000000000000000000000000110100000001000000000000000100000000111100000000000000010000000000000000000100001101000000001101000100000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000001111000100001111000000000000000111111111000000000000000000010000000000010000000011110000",
		"00000000000000010000111100000000000000000000000000000000111000010000000000000000000000001111000000000000000000000000000000011100000011100000000000000000000100000000000000000000000000000000000000000000111100000001000000000000000000000001000000000000000100010000000011110000000000001110000000001111000000011111001000000000000000010000111100001111000011110000000000000000000000000000000000000000000000000000111100000000000000000000000100000000000000000000000011110000111100001111000100000000000000010000000100000000",
		"00000000000000000000111100000000000000000000000000010000111100000000000000010000000100000000000000000000111100000000000000011011000011010000000100000000000100000000000000000000000000000000000000000000000000000001000000000000000000000001111100000000000100010000000011100000000000001110000000001111000000000000001011110000000000000000000000000000000011100000000100000000000000010001111100000000111100000000000000000000000000000000000100000000000000000000000000000000111000000000000000000000000000000000000011110000",
		"00010000000000001111000000000000000000001111000000000000111100001111000000000000000000010000000000000000000000000000000000001100000011100000000000000000000100000000000000000001000000001111000100000000000000000000000000000000000000000001000011110000001000010000000011110000000000001110000000010000000000000000001011010000111100001111000000001111000011110000000000001111000000100001000000000000000000000000000000000000000000000001000000010000000000000000000100000000000000000000000100000000000000000000111011110000",
		"00010000000100000000111100000000000000000000000000010000000000000000000100000000000000000000000000000001000000000000000100001101000011100000000000000001000100000000000000010000000000000000000000000000000000001111000000000000111100000001000000000000000000000000000000000000000000010000111000010000000000000001000111010001000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000111100000000000000000000000000000000000100000000000000001111000000000000000000000000111000000000",
		"00010000000100000000111100000000000100000000111100010000000000010000000000000000000000000000111111100001000000000000000000001110000011110000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000010000111100000000111100000000000000000000000000000000111100000000000000000000001011110000000000000000000000000000000000010000000000000000000000010000000000000000000011110000000100100000000000000000000000000000000000000000001000000000000000001111000000000000000100000000000000000000",
		"00000000000100000000111100000000000000000000111100010000000000100000000000010001000000000000000000000001000100000001000000000000000000000001000000000001000000000000000000001111000000011111000000000000000000000000000000010000000000000000000000000000111100000000000000010000000000000000111100000001000000010000000100000000000000000000000000001111000100100000000000000000000000000000000000000000000111110000000000010000000000000000000000010000000000000000000100000001111100000000000000000000000000000000000000000000",
		"00001111000100000000000000000000000100000000000000000000000000010000000000000001000000010001000000110000000000000010000000000000000000000000000000000000000000000001000000010000000000010000000000000000000000000000000000000000000100010000000000000000111100000000111100000000000000000000000000000000000000000000000011110000000000010000000100000000000000010000000000000000000000010000000000000000000000000000000000000000111100000000000000000000000000000000000100000000000000010000000000001111000000000000000000000000",
		"11110000000000000001000000000000000100010001000000000000111100000000000000000001000000010000000100110000000000000001000000000000111100000000000000000000000000000001000000010000000000010000000000000000000000000000000000010000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000010000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000011110000",
		"00000000000000000001000000001111000100000010000100000001111000000000000100000000000000000001000000010000000000000000111100000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000100000000000100010000000000000000000000001111000000000000000000000000000000000001000100001111000000000000000000000000000000000000000000010000000000001111000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000",
		"00000000000000000000000000000000000100000000000100000000111100000000000100000001000000000000000000000000000000000000000000000001000000000000000000000000000111110001000000010000000000000001000000000000000000010000000000011111000000001111000000000000000000000000000000000001000000001111000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000011111000000011111000000000001000000001111000000010000000000000000000000000000000000000000000000010000000011110000000100001110000011110000",
		"00000000111100000000000000000000000000000000000000001101000000000000000100000001000000000001000000000000000000000000000000000001000000000000000000000000000100000001000000000000000000000000000000001111000000000001000000000000000000000000000000000000000000000000000100000001000100000000000000000000000000000000000000000000000000010000000100010000000000010000000000000000000000011111000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011110000",
		"00001111000000000000000000001111000100001111000000011101000000000000000000000000000000000000000000000000000000000000000100000000000011110000000000000000000100000000000100010000000000000001000000001111000000000000000000000000000100000001000000000000000000000000000000000000000100001111000000000000000000000000000000000000000100010000000100010000000000001111000000000000000000011111111111110000000000000010000000011111000000000000000000000000000000001111000000000000000000010000000000000000000000001111000000000000",
		"00000000000000000000000000001111000000001111000000001110000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000001111000100000000000100000000000000000001000000001111000000000000111100000000000100000010111100000000000000000000000000000000001000001111000000000000000000000001000000000000000100011111000000010000000000011111000100000000000000000000000000000000000000000001000000011111000000010000000000001111111100000000000000000000000000000000000000000000000000010000000100000000",
		"00000000000000000000111100000000001000001111000000001111000000010000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000100000001000100000000000000000000000011111110111100001111000000000000000100000000000000001111000000000000000011110000001000001111000000000001000011110000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000011110000000100000000000001110000000000000000000000000000000000000000000000000000000000010000000000001",
		"11110000000000000000000000001111000100000000000000000000000000010000000000000010000000000000111100000001111100000000000000000001000000000000000000000010000111110000000000000000000000000000000000000000111100001111000000000000001000000001111100000000000011110000000000000000000100000000000000000000000011101111000000010001000000100001000000000000000000000000000011110000000000010000000011110000111111110001111100011111000000100000001000000000000000001110000011110000000000000000000011110000000000000001000000000001",
		"00000000000000000000000000001111000000000000000000000000000000000000000000000010000000000000000000010000000100010000000000000000000000000000000000000001000000000000111100011111000000000000000000010001000000000000000100001111000000000000000000000000000100000000000000010000000011110000000011110000111100000001000000010000000000000010000000000000111100000000000100000000000000011110000011110000000011110001000000000000000000100000001011110000000011111111111100001111111111111110000000000000000000000000000000000001",
		"00000000000000000000000000010001000000001111000100000000000000000000000000000001000100000000111100010001000000010010111100000000111100000000111000001111000000001110111011111111000011110000000100000000000100011111000011110000000000000000000100000000000000000001000000010000000000000001000000000001000000000001000000100001111100000001001011100000111000000001000000010000000000001110001011110000000000000001000100000000000100100000000011110000000011100000000000001111111100001110000011100000111100000000111000010000",
		"00001111000000000000000000000000000000000000111100000000000000000000000000000000000000000010000000001111000000000000000000000000000000000000111000000000000000001111000000000000111100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000010000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00001111000000000000111100000000000100011111000000000000000000000000000111110000000011110000000000000000000100010001000100000001000000000000000000000000000000000000000000001111000000010000000000000000000000000000111100000000000000001111000000000000000000000001000000010001000000000000000000000000111100010001000000000001000000010001000000000000000000000000000100010000000000000000000000000000111100000001000100000000000011110000000100000000000000000001000000001111000000010000000011110001000000010000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000100000000111000011110000111100000111100010000111100010000000100000001000000001111000011110000000000000001000000000001000000000000000000000000000111110000000111110001111100000000000000000000000000010000111100000000000000010000000000000000000011101111001011110010000000000000111100010001000000001110000100000000000000100000000000010000111100001111000100010000000111110001111100000001000011110000000000000000000100000000000000000000111100000000000000000001000000000000000000000000000100010000000100000000",
		"00001111000100000000000000011111000100001111111100000000111100010000000000000001000011110000000011111110000100000000000000000000111100000000000000000000001000000000000011110000000000000000000000000000000000000000111000010000000000010000000000000000000011111111000100000010000000000000000000000001000000001111000000000000000000010000000000000000000000000000000000010000000000000000111100000000000000000001000000001111000100000000000111111111111100001111000100000000000000000000000000010000000000010000000100000000",
		"11110000111100000000000000001111000100001111000000001111111100010000000100000000000000000000000000000000000000000001000000000001000011110000111000001110000000000000000000000000000000000001000000001111000000000000111000010000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000011110000000000000000000100000000000000000000000000000000000000001111000000000000111100000000000000000000000000011111000111101110000000111101000011110010000000000000000000001111000000000000000000000001",
		"11110000111100000000000000000001000011110000000011110000000000000000000000000000000111110000000000010000000000010000000000000000000011100000000000000000000011110000000011110000000011110001000000010000000000000000000000000000000000000000000000010000000000001111111100000000000000000000000000000000000000000000000000000001000000000001000000010000000000000000000000010000111111110000000111110000000011110000000000000000000000001111000100001110111100011111000100000000000000000000000000001111000011110000000000000000",
		"00000000111100000000000000001111000100000000000000000000000000000000000000000000000000001111000100000000000000000001000000000000000011110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000001111000011110000000100000000000000000001000000001111000000000000000100000010000000000000000000000000000000000000000000000001000000000000000011110001000000000000000000000000111111110000000000010000000100000000000000010000000000000000111100000001000100000000",
		"00000000000000000000000000000000001000000000111100000000000000010000000011110000000000001111000000000000111100000001000100000000000011100001000000000000000000000000000100000000000000000001000000000000111000000000000000010000000000000000111100001111000000001111000011110001000100011111000000001111000000000000000011110000000000000001000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000001111000000000000000000010000000111110000000000010000000000000000000000010000000111111111",
		"00000000000000000000000000000000001000000000000000000000111100000000000000000000000000011111000000000000000000000001000000000001000011010000000000000000000000000000000011110000000000000000000000010000111000000000000000000000000000000000000000000000000100010000000000000000000000001110000000001101000000000000000111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000011111111",
		"00000000000000000000000011110000000100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000100000000000000000000000111110000000000000001000000000000000000000000000000000000000000000000000000000000000100010001111111110000000000001110000000001110000000000000000111100000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100000000000000000000111100000000000100000000000000000000000111100000",
		"00000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000001000000010000000000000000000011110001000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000100010000000011110000000000001111000000011110000000000001001011110001000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000000000000100000000000000000000000100000000111100001111000000000000000000000000000011100000",
		"00010000000000001111000000000000001000001111000000000000000000010000000000000000000000000001000011110001000000000000000000000000000000000001000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111100011110000000000000000111010000000000000000000000000000000000000000000011110000000000000001000000001111000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000011110000",
		"00000000000000001111000000000000000100001111000000000000000000000000000000000000000000010000000011110001000000000000000000000000000000000001000000000000000100000000000000000000000000000000111100000000000000000000000000010000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000111010000000000000000000000000000000000000000000011110000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001111000000000000000000000000111100000000",
		"00010000000000000000000000001111001011110000000000010000000000010000000000000000000000000000000011110001000000000000000000000000000000000001000000000000000100000000000000000000000000000000111100000000000000000000000000000000000000010000000000000000111100000000000000000000000000000000111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100010000000000000000000000000000000000000000001000000000111100001111000000000000000000000000111100000000",
		"00010000000100010000000000001111000100001111111100000000000000101111000000000001000000000000000000000000000000000001000000000000000000000000000000000001000000000001000000000000000000000000111100010000000000000000000000000000000100010000000000000000000000010000000000000000000000000000111000000000000000000000000011110000000100010000000000000000000100000000000000000000000000010000000000000000000000000001000100010000000000000000000000000000000000000000000100000000111100000000000000000000000000000000000000000000",
		"00000000000100000000000000001111000100001111000000000000000000010000000000000001000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000010000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000100010000000000000000000000010000000000000000000000010000000000000000000000000010000100001111000000000000000000000000000000000000000100000000000000000000000000000000000000000000111111100000",
		"00000000000100010000000000000000000100000000000100000000000000000000000000000001000000000000000000100000000000000001000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000100010000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000111111110000",
		"00000000000000000000000000001111000100000001000000000000111000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000001000100010000000100000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000010000000000000000000000010001000000000000000000010000000000000000000000000000000000000000000000000001000000000000000100000000000011100000",
		"00000000000000010000000000000000000111110000000000001110110100000000000100000001000000000000000000001111000000000000000000000000000000000000000000000001000100000001000000000000000000000000000000001111000000010000000000000000000000010000000000000000000000010000000000000001000000001111000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000010000111100000000000000001110000011100000",
		"00001111000000000000000100000000000100000000000000001100111100000000000000000000000000000000000000001111000000000000000000000000000011110000111100000000000000000001000000010000000000000001000100001111000000000000000000000000000000010000000000000000000000000000000000000000000100001111000000000000000000000000000000000000000000010000000000000000000000001111000000000000000000010000000000000000000000000001000000000000000000010000000000000000000000001111000000000000000000010000000000000000000000001110111111100000",
		"00001111000000000000000000001111001000000000000000001101000000000000000000000001000000000000000000011111000000000001000011110001000011110000000000000000001000000000000000000000000100000010000011111111000000000000111100000000000000010000000000000000000000000001000000000000001000000000000000000000000000000000111100000000000000010000000100000000000000000000000100000000000000010000000011110000000000000001000000001111000000000000000000000000000000001111000011110000000000000000000011110000000000000000000011100000",
		"11110000000000000000000000001111000000001111000000001110000100000000000011110000000000000001000000000000000000000000000000000000000000000000111100000000000100000000000000010000000100000001000100001111000000000000000000000000000000000010000000001111000011110000000000000000001000000000000000000000000011110000000000000000000000010000000000000000000000011111000000000000000000000000000111100000000000000000000000000000000000000000000000001111000000011111000000000000000000010000000011111111000000000001000011110000",
		"00000000000000000000000000001111000000001111000000001111000000010000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000100000000000000000001000100000001000000000000000000001111111100000000000100000001000000000000000111111111000100000001000100000000000000000001000111111111111100000000000000010000000000000000000000001111000000000001000000000000000011110000000000000001000000010000000000000000000100011110000000011111000000000000000000000000000011110000000000000001000011110000",
		"00000000000011110000000000000000000100001111000000001111000000000000000000000001000000000000000000000000000000000001000000000000000000001111000000000000000000000000000000000001000000000000000000000000111100001110000000010000001000010000000000000000000100000000000000000000000100010000000000000000000111100000000000010001000000010001000000000000000000000000000011110000000000000000000011110000000000000001000000010000000000011111000100000000111100011111000000000000000011111111000011100000000000000000000000000000",
		"11110000000000000000111100010001000000001111000100000000000011110000000100010001000100000000000000100000000100010000000000000000111100001110111100000001000000010000111100011111000000000000000000000000000000011111000100000000000000100000000000000001000100000000111100010000000000000001000000000000000011110001000000000010111100000010000000010000111000000000000000000000000000001111000111110000000011110001000011110000000100101111001000000000111100001110000000001110111100001111111011101111000000001111000000000001",
		"00001111000000001111111100000001000000101110000100010000000000001110000100000000000100010000000000010000000011110001000000000000111000010000111100001111000000010000111100000000000000000001000111110000001000100000000011110000000000010000000000000000000000000001000000001111000000000001000100010000000011110000000000000001111100000000000111100000111000000000111100100001000000010000000000000000111100000001000000000000000100100000000100000000000000000000000000001111111000001111000111111111000000000000111100000000",
		"00010000000000000001111100000000000000000000111100100001111100001111000100000000000000000001000000001111001000011111000000011111000000000000000111111101001000010000111000000001000100001111000000010000000100001110111100011111111100010001000000000000001000011111001011110010111100011110111100100000000100000000111111110010000000001111000000011111000000001111000000100000000100000001111100010000000011110000000000001111000000000000000011100000111000000010000000010000000111100000001000001111001100010000000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00001111000000010000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000011110000000000000001000000000001000000000001000000001111000000000000000000000000000000000001000000000000000000000000000000001111000000000000000000000000000000000000000000000000000011110000000000000000000000000001000000000000000000000000000000000001000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000000000000111100000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000011110000000000000000000000000000000000000000111100000000000000000000000000001111",
		"00000000000000000000111100010000000000000000111000000000000000000000000000000000000000000000000011100000000000000000111100000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000100000000000000000000000000000000001011110001000000000000000000000000000100001111000000000000000000010000000000000000111100000000000000010000000100000000000000000000000000000000000011110001000100000000000000000000111100000000000000000000000011110000000000000000000100000000000000001111",
		"00001111000000000001000000001111000100011111111000010000111100000000000011110000001100000000000011111111000011110001000000000000111000000000001000000000001000001111000011110001000000000000000011110001000000000000111000011111000100010000000000000001000000000000000011110000000000000000111100000000000100001110000000001111000000000000000100000000000000000000000000000000111100000000000000001111000000000001111100000000000000010000000000000000111100010000000100000000000000000000000100000000000100000000000000000000",
		"00001111000000011111000000011111000000010000111100000000000100000000000000000000000100001111000000000000000011110001000000000001000011110000000000000000000011110000000111111111000011110000000000000000000000000000110100010000000000000000111100000000000000000000000000001111000000010000000000000000000000001111000000000000000000010001000111110000000000000000000000000000000011110000000000011111110100000000000100000000000000001111000011111111000000101110000000000001000000001111000011110000000000010000000000000001",
		"00001111000000000000000000001111000100001111000011101111000000000000000000000000000011110000000100001111000000000000000100000001000011100000000000000001000000000000000000001110000000000000000000010000111100000000000000010000000000011111000000001111000000001111000011110000000000000000111100011111000000001111111100000010000000000011000100000000000011110001001000000000111100000000000000000000111000000001111111110000000000001111000100001111000000101110000111110000000000101111000011111111000100010000000100000000",
		"00000000000011110000000000000000000100001111000011111111000000000000000000000000000011110000000100000000000000010000000100000001000011110000000000000000111100000000000111111111000100000000000000010001000000000000111100000000111100001111000000000000000000001111000011100001000100011111000000000000000000000000000000000000000000000010000000000000000000000001000111110000000000000000000000000000111111110010000000000000000000000000000011110000111100101111000100000000000000001111000000000000000000000001000100000000",
		"00001111000000000000000000000000000100000000000000000000000100000000000000000000000011110000000000000000000000000000000000000000000011110000000100000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000001111000000010000000011110000000100100000000000001111000100000000000000000000000100000000000000000000000000000000000011110000000000000000000000000000000000000001000011110000111100000000000000001111000000101111000100000000000000000000000000000000000000000001000000000000",
		"00000000000011110000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000111100000000000011110000000100000000111000010000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000001111000000000001000000000000000000000000000011110000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000001111000000000000000000000000000011110000",
		"00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000010000000000000000111100000000000000010000000000000000000000010000000000000000000000010000000000001110000011110000000011010000000000010000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000001111000100000000000000000000000011110000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000000000000000000010000000000000000000000000000000000000000011110000000000000001111100010000111100000000000000010000000000000000000000000000000100000000000000000000000000010000000100001111000000000000000011100000000000001111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000001111000000000000000000000001000111110000",
		"00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000001000100000000000000000000000000000000000000000001111100010000111100000000000000010000000000000000000000000000000000000000000000000000000000000000000000001111000000010000000011010000000000001111000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000001000000010001111100000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000011100000000000001111000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000010000000000000000000000000001",
		"00000000000000000000000000001111000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000100000000000000000000000000000001111000000000000000000000000100010000000100000000000000000000000000010000000000000000000000000000000000010000000000000000000011110000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000001000000000000011110001000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001111000000000000000000000000100010000000100000000111100000001000000000001000000000000000000000000111100000000000000000000000000000000000100000000000000000000000000000000000011110000000000000000000000000000000000010010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000",
		"00000000000100000000000000000000000100001111000000000000000000010000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000100000000000000010000111100010000000000000000000100000000000000000000111100010000000000000000000000001111000000000000000000000000000000010001000011110000000000000000000000000000000000000001000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000111011110000",
		"00000000000000000000000000000000000100000000000100000000000000010000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111100010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000010001000000000000000000000000000000000000000000000000000000000000000000001111111111100000",
		"00000000000000000000000100000000000100000001000000001111111100000000000000000001000000000000000000010000000000000001000000000000000000000000000000000000000000000001000000010000000000000000111100000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000111100000000000100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000001111000000010000000000000000000000001111000011110000",
		"00000000000000000000000000000000000000000000000000001101111000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000100010000000011110000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000010000000000010000000000000000000000001111000100000000000000000000000000001111111111100000",
		"00000000000000000000000000000000000000011111000000001110000000000000000000000000000000000001000100001111000000000001000000000000000011110000000000000000000100000001000000010000000000010000000000001111000000001111000000000000000000010000000000000000000011110000000000000000000100001111000000000000000000000000000000000000000000010000000000000000000000001111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000011110000",
		"00001111000000000000000000000000000100001111000000001110000000000000000000000000000000000001000000000000000000000001000000000001000000000000111000000000000000000000000000001111000000000010000000000000000000001111000000000000000000010001000111110000000011110000000000000000000100000000000000000000000000000000111100010000000000010001000000000000000000001111000000000000000000010000000000000000111111110000000100000001000100000000000000001111000000001111000000000000000000010000000011110000000000000000000000000000",
		"11110000000000000000000000010000000000010000000000001110000000000000000011110000000000000010000000000000111100010000000100000000000011110000111100000000000000000000111100000000000100000001000000001111000000011111000000000000000100000001000100001111000011100000000000010001000100000000000000000000000000000000000000000000000000010001000000010000000000011111000100000000000000010000000011110000000000000000000000000000000000000000000000001110000000000000000000000000000000010000000011110000000000000000000000000000",
		"00000000000011100000000000000000000000000000000000000000111100000001000000010000000000000000111100000000000000000000000000010000000011110000000100000000000011110001000000000001000000000001000100000000000000001110000000000000001000010001000000000001000011110000000000000001000100000000000000000000000111111111000000000000000000010001000000000000000000010000000000000001000100000000000011110000000011110000111100000000000000000000000000001110000000011111000000000000000000000000000011100000000000000001000011110000",
		"00000000000011110000111100000000000100000000000000000000000000000001001000010010000100010000111100000000000000000000000000000000111100000000000000000001000000000001000000000000000111110001000011110001000000001111000000010000001100100000000000000000000011110001111100000000001000010000000000000000000111110000000000000001000000000001000100000000111100000000000011110001000100001111000111100000111100000001000000000000000000100000001000000000000000011111000000001111000011100000000011100000000000000000111111110000",
		"11110000000011100000000000000000000000000000000100000000000000000001000100100000001000000001000000010000000011110001000011110000000000001111111100000000000000001110000000010000000011110001001000000001000000010000000011110000001000010000000000010001000011110000111000000000000100010001000000001111000011110000000000000000111100000010000100010000111100000000000011110001000000011110001011100000111111110001000000000000000000010000001000000000111100011111000100001101000011110000111011100000000011110000000000000000",
		"00001111000100001111000000000001000000010000000100000000000000000000000100010000000100000001000000010000000011100001000011100000111100000000000000000000000000000000000000010000000111110001000011111111000000010000000000000000000100010000000000011111000011100001111100001111000100000001000000001111000000000000000000000000111100010001000000000000111000010001111100000001000000010000000000001111111100000011000000000000000100010000000100000000111100000000000000001110111100001111000000000000000000000000111100000000",
		"00100000000000001111000000000000111100001111000000000001000000001111000000001111111100000000000000000000000000001111000000000000000000000000001000001110000111110000111100000000000000000001000000001111000000010000000000000000111100010000000000001111000000000000111111110001000111110000111100010001000000010000000000000000000000000000111100000000111100000000000000000000000000000000000011110000000000000000000000001111000011110000000000000000111100000001000000000000000000000000000111111111000100000000111100000001",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000111100000000000000001111000000010001111100010000000000000000000000000000000000000000000011110001000000000000000000000001000000000000000000000000000100000000000000000001000000000000111100010000000000000000000000000000000000001111000011111111000000000001000000001111000000000000000000010000000100001111000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000100010000000000000000000000011111111111110000",
		"00000000111100000000000000000000000000001111111100010000111000000000000000000001000000000000110100000000000011010010111111110001110100010001000100000000001000000000000111110000000011110000000011110001000000000000000000010000000100000000000000000000111100001111000011110000000000001111000011110000111100001110001000001111000000001111000000000000111100000000000000000001000000000000000000001111000000000000000000100000000000011111111100011111111100000000000111110001000000000000000000000000000000001111000000000000",
		"00100000111000001110000000011110000000011111111100011111000000000000111100000000000000000000000011110001111011100010000000000010111000000001000100000000000000000000000011110000111100000000111100000000111100000000111000010000000100010000000000000000111100001110000011101111000000001110000000000000000000001110000000011111000000010000000000000000111100000000000000000000000000000000000000000000110100000000000000000000000000000000000000001111111100100000000100000000111100000000000011110000000000010000111100000000",
		"00000000111100001111000000001110000000000000000000000000000011110000000000000000000011110000000100000000111100000001000000000010111100000001000000000010000000000000000011110000111100000000111100000000111000010000111100000000000000011111000000001111000000011111111100000000000000001111000000010000000000011111000100000000000100000010000000000000000000000000000000000001111100000000000000000000111000000000000000000000000000000000000100000000111100000000000011110000000000011111000000001111000000010000000000000000",
		"11111111000000000000000000000000000000000000000000001111000000000000000000000000000000000000000100000000000000000000000100010001000000000000000100000001000000010000000011111111000000010000000000000000111000000001111100000001000000000000000000010000000000001111000000000000000000010000000000010000000000000000000000000000000100000001000000000000000000000000000000000000000011110001111100010001000000000001000011110000000000000000000011111111111100000000000000000000000000011111000000001111000000000000000000000000",
		"00000000000000000000000000000001000000000000000000000000000000000000000000000000111000000000000100000001000000010000000000000000000000010000000000000000000000001111000000000000000100010001111100000000110100010000111100000000000000000000000000010000000000001111000000000000000000001111000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000111000000001000000000010111100000000000000000000111100000000000000011111000000000000000000000000000000000000111100000000000011111111",
		"11100000000011110001000000000000000000001111000000000000000000000000000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000001111000000000000000100010001111100000000000000000000111100000000000100000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000011110000000011110000000000000000000000000000000000000000111000000000000000000000000000000000000000011111000000000001000000000000000100000000111100000000000011110000",
		"00000000000000000000000000000000000000000000000000000000000011110000000100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111100000000000000000000111000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000011110000000000000000000000000000000000010000000000000001000000000000000000000000000000000001000000100000000000000000000000000000000111110000000000000000000111110000",
		"11110000000000000000000000000000000000000000000000000000000000000000000100000000000000000000111100000000000000000000000000000001000000000000000000000000000000000000000011110000000100000000000000000000000000000000111100000000000000001111000000000000000011110000000000000000000000000000000100000000000000000000000011100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000111100000000000000000000",
		"00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000010000000000000000000000000000000000000000000000001001000000000111100000000000000000000000000000000000000010000000000000001000000000000000000000000000000010000000100001111000000000000000011110000001000001111000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000100000001000000000001000000000000111100000000000000000000",
		"00000000000000000000000000001111000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000001000000000000000100000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000100000000000011110000000000001111000000000000000000000000000000000000000000000001000000000000000000000000000000001111000000000001000000000000000000010000000000000000000000000000000000000000000000000000000011110000",
		"00000000000000000000000000000000000000000001000011110000000000000000000000010000111100000000000000000000000000000000000000000001000000000000000000000001000000000000000000000001000100000000111100000000000000000000000000000000000100000000111100010001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000011110000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000",
		"00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000100000000111100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000011110000000000000000000100000001000000000001000000000000111100000000000000000000000100000000000000010000111100000000000000000001000000000000000000000000111100000000000000010000000000010000000000000000000000000000000000000001000011110000000000000000000000000000111100000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111100000000",
		"00000000000000000000000000001111000100000000000100001110000000000000000100000000000000000000000000010000000000000001000100000000000000000000000000000001000100000000000000000001000100000001111100000000000000000000000000000001000000010000000000000000000000000001000000000000000100000000111100001111000100000000000100000000000000000000000000000000000000000000000011110000000000000001000000000000000000000000000000000000000000000000000000000001000000001111000000000000000100000000000000000000000000001111111100000000",
		"11110000000000000000000000001111000100001111000000001101111000000000001000000000000000000000000000010000000000000000000000000000000100000000111100000001000100000001111100000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000001111000100000000111100000000000000000000000100001111000000000001000000000000000000000000000011100000000000010000000000000000000000000000000000000000000000000000000100000000000100001111000011111111000100000000000000000000111100001111111111111111",
		"11110000000000000000000100000000000000000000000000001110110100000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000001000000010000000000000001001000000000000100000000000000000000000000000001000100001111111100000000000000001111000000000000111100000001000000000000000111110000000011110000000100000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000100010000000000000000000000001111000011101111",
		"11110000000000000000000000000000000000010000000000001110111011110000000000000000000000000000000100010000000000000000000000000000000011110000000000000000000000000000000000000000000100000000000000000000000000010000000000000001000100010000001011101111000000000000000000010000000100001111000000000000000000001111000000000000111100000001000000000000000000001111000011110000000000010001000000000000000000000000001011110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000011110000000000000000000100000000000000001111111100000000000000000001000100000000000000000000000000000010000000000000000011110000000000000001000100000000000000010000000000000001000000010000000000001111000000000000000100000000000111110000000000000001000000010000000000011111000000000000000000001111000000000000000000100001000000000000000000011111000100000000000000010000000100001111111100000000000000000001000100000001000000000000000000001111000011110000000000000000000011110000000000000000000011110001",
		"00000000000011110000000000000001000100010000000000001111000000000001000000000000000011110010000000000000111100000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000001100000000000100000000000011110000000000000001000000010000000000000000000011110000000011110000111000010001000000000000000000011111000100000000000000001111000000000000000000000000000000000001000000000000000000001111000000000000000000000000000000000000000011100000000000001111000011111111",
		"00000000000011100000000000000000000100000000000011110000000100000001001000000000000100000000111100000000111100000001000000000000000011110000000000000001000000000000000100010000000011110000000000000000001000001111000000001111001000010001000100000001000000000000000000000000000100010000000000010000000011110000000000010000000000000000001000000001000000000000000111110000000000001111000000000000111011110000111100000000000000101110111100001111000000000000000000000000000000000001000011100001000011110000000011111111",
		"00000000000011100000000000000000000100000000000000000000000000000001001000010001000100001111111100000000111100000010000011110000000011110000000000000001000011111110000000000000000000000001000100000000001000000000000000000000001000010010000000010000111100000001111000001111001000010000000000101111000011111111000000000000000000000000000100000001000000000000000011110010000000000000000111110000111100000001000000000000000000101111000100010000000000011110001000001110000111110010000011100000000000000001111111101111",
		"11100001000000000001000000000000000000000000000100000000000000000001000100100000001000000000111000000001111100000001111011110000000000000000000000000000000000001110000000000000000011100001000100000000001000010000000100000000000100010000000100010000111100000001111100001111000000000000000000000000000000000001000000000000000000000010000011110000111000000000000011100001000100001111000111100000111111110001000011110001000100001111001011110000111100001110000100000000111100000001111011110000000000000000000000000000",
		"00000000000000000000000000000001000000010000000100000000000000000000000100010000000100000000000000010000000011110000000011110000000000010000111100001111000000000000000000000000000100000001000111111111000000000000000000000000000000010000000100011111111111110000111111111111000000000000000000011111000000000000000000000000000000010000000000000000111100000000000000000000000000000000000011110000000000000010000000000000000000010000000000000000111100001111000100000000000011110000000000000000000011110000111111100000",
		"00010000000000011111111100010000111100001111000000001111000000001111000100000000111100000000000000000000000011110000000011110000000000000000000000000000000011110000000000000000000000010000000011111111111100010000000000000000111100011111000011110000000100000001000000010000000011100001000000010000111000010001000000000001000000000001111111110000111000000000000000010000000000000000000100001111000000000000000100000000000000000001000100000000111100000000000000001111000000000000000011110000000100000000111100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00011111000100001111000000010000000000000000000100010000000100001111000000000000000000000000000100000000000100001111000000000000000100000000000011110000000000000000111100001111000011110000000011110000000000000000000000000000000011110000000000000000000000000000000000000000111100000001000000000000000011110001000011111111000000001111000000010000000100000000111100001111000000000000000000010001000100001111000011110001000111110000000011111111000000000000000000000000111100000000000000000000000000010000000000000000",
		"00000001000100010000000000100000111111110000000000010000000000000001000000010000111100001111000000010000001011110000000000000001000000000001000000000001000000000000000011101111000011110000000000000000000000000001000000010001000000000000000000000000111000001111000000000000000000000001000000000000000000011111001000011111000000000000000000000000000000000000000000000000000000001111000000010000000100000000000000000001000011110000000000001111000100000000000100000000000100000001111100000000000000000000000000000000",
		"00000001000000000000000000100000111011110001000000000001000000000000111100010000000000000000000000010001111100010000000011110010000000010001000000000001000000010000000011100000111011101111000000000010111111110001111000010001000000100001000100000010111100010000000000000000000000010000111100000011000000100000001000010000000100000000111100000000111100000000111111110000000000000000111100000010000000000000111100000001000111101111000000001111000011110000001000000000000000010000111000000001111100000000111000001111",
		"00000001000100001111000000000000111100000000000100000010001011100000111000011111000000000000000100100000111000000000000000000001000000010001000000000001000000010000000011101111111111110000111111110001111000000001111100000001000000000000000100000001000000010000000000000000000000010000000000000000000000000000001000000000000000000000111100000000111100000000000000000000111100000000000000000000000000001111000011110000111100001111000000000000000000000001000100000000000100001111111100000000000000000000111100001111",
		"00000000000100010000000000000000000011110000000000001111000100000000000000010000111100000000000000000001000000000000000000000001000100010000000100000001000000010000000000000000000000010000111100000001110100000010000000010000000000000001000000010000000000000000111100000000000000000000000000000000000000000000000000010000000100000001000000000000000000001111000011110000000011100000111100010000000000000000000000000000000011110000000011100000000011110001000100000000000100000000000000000000000000000000000011110000",
		"11110001000000010000000000000001000000000000000000000000000100000001000000010001111100000000000000000001000000010000000000000001000000010000000000000001111100000000000011110000000000000000111100000001110000000010111100010000000000010001000000010001000000000000000000000000000000000000000000000000000000000001000100000000000000000001000000000000000000001111000011100000000011110000111100000000000000000000111100001111000011111111000000000000000000000000000100000000000000000000000000000000111111110000000000000000",
		"11000000000100000000000000000001111100000000000000000000000100000001000000010000111100000000000000000001000000010000111100000000000000000000000000000000111100000000000000000000000100000001111000000000111000000001111000000000000000000000000000010000000000001111000000000000000011110000000000000000000000000000000100100000000000000001000000000000000000000000111111110000000000000000000000000000111111110000111100000000000000001111000000000000000000000000000000000000000000000000000000000000111111110001000011111111",
		"11010000000000000000000000000001000000000000000000010000000011110000000000010000000000000000000000000000000000010000000000010001000000000000000000000000000000000000000000000000001000000001111000000000000000010001111000001111000100000000000000100000000000001111000000000001000111110000000000000000000000000000000000011111000000000001000100010000000100000000000000000000000000000001000000010000111100000001111100000000000000000000000000000000000000011111000011110000000000000000000111110000000011110000000000000000",
		"11100000000000000000000000000001000000000000000000000000000000000000111100010000000000000000000000000000000000100000000000000010000000000000000000000001000000000000000000000000000000000000111100000000000000000001111100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001111000000000001000000000000000000000000000000000000111100000000000000000000000011110000000000000000000000000001000000000000000000000000000011110000000100010001000011110000111100000000000100001111",
		"00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000111100000000000000010000000000000001000100000000000000000001000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000010000000000000000111100000000000000000000111100000000000100001111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000100100000000000000000000100010001000000000000111100000000000100001111",
		"00000000000000000000000000000000000100000000000000000001000000010000000100000000000000000000111100000000000000000000000000010001000000000000000000000001000000000000000000010001001000000010000000000000000000000000000000000000000000000000000000000000000000001111111111110000000100000000000000010000000100000000000000000000000100000000000000010000000100000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000010000000000001111111000000001000100000000",
		"00000001000000000000000000001111000000000000000000000000000000000000000100101111111100000000000000000000000000000000000000000000000100000000000000000010000000000000000000000001000100000000000000000000000000000001000000000000000000000000000000010000000000000000111111110000000000000000000000000000000100000000000000010000000000000000000000010000000100000000000000000001000000000001000000000000000000000001000000010000000000000000000000000000000100000000000000000000000100000000000011110000111100000001000000010000",
		"00010001000000010000000000000000000000000000000000000000000000000000000100100000111100000000000000000000000011110000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000100010001000000000000000000010000000000000000000000000000111111110000000000000000000000000000000000001111000000010000000000000000000000000000000000000000000000000000000000010000000100000000000000010000000000010000000011110000000100000000000000010000000000000000000000010000000000000000111100010000000000010000",
		"00010001000000000000000000001111000100000000000100000000000100000000000100000000000000000000000000010000000000000000000000000000000000000000000000000001000100000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000010001000011110000000000000000000000000000000000000000000100000000000000000000000000000000111100000001",
		"00000010000000000000000000000000000100000000000100001110111000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000111100010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000111110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011110000000000000000000000000000000000000000000000010000000000000000000000001111111100000000",
		"00000001000000010000000000010000000100001110000100001110110100000001000100000001111100000000000000010000000000000001111100000000000000000000111100000000000100000001000000000000000000000000000000000000111100000000000000010000000000100000000000000000000000000000000000000000000100000000111100000000000100000000000100001111000000010000000000000000000000000000111100000000000000010000000000000000000000000000000000000000000111110000001000001111000000000000001000001111000000000000000000000001111100001111000000000000",
		"00000000000000000000000011111111000000001110000000001110110100000000000100000000000000000000000000000000000011100001000000001111000000000000000000000000000000000001000000010000000100010000000100000000000000011111111100000000000100010000000100000000000000000000111100000001000000001111111100000000000000000000000100001111000000000000000000000000000000001111000011100000000000000001000000001111000000000000000100000000000000000000000000001111000000000000000111110000000000000000000000000000111100001111000000000000",
		"00000001000011110000000011100000000000010000000000001101110100000000000000010000000000000000000000000000000000000001000000001111000000001111000100000001000000000000000000010000000000000000001000000000000100000000000000001111000000010000000100000000000000000000111100000000000000001111000000000000000000000000000000000000111100000010000011100000000000010000000011110001000000010010000100000000000000000000000100000000000000000001111100000000000000000000000100001111000000000000000000000000111100001110111000000000",
		"00000001000011110000000000000000000000000000000011111111000000000001000000010001000000000000000000000000000000000010000000000000000000000000000100000001000000000000000000000000000100000000000000000000000000000000000000000000000100000000000100000000000000000000000100000000000000001111000000000000000011100000000000001111000000000001000111110000000000000000000100000001000100000000000100000000000000001111000000000000000000000001000000000000000111111111000000000001000000000001111100000000111100001111111111110001",
		"00000001000011110000000000000001000000000001000000001110000000000010000100000000000000000010111100001111000000000001111100000000111100100000000100000010000000000000000000000000000000000000000000000000000000000000000000001111000000000000001000000000111100000000000000000001000100000000000100000000111011110000000000000000111100000010000011110000000000010000000100010000001000001111000000010000000100000000000000000000000000000000000100000000000000000000000011110000000000000010111111110000000011111111111000001111",
		"00010001000000000001000000000001000011110000000111111111000000000010000000010000000000010000111100100000000000000001111100000001000000011111000000000010000000000000000000000000000000000000000000000000000000000000000100001111000100000000000100010001000011110000111100000000000000000000000100000000111000000001000100001111000011110000000000000000000000000000000000000000000000001110000100001111000000000000000011110000000000100000000000000000000011111111000000000000000111110010111111100000000011101111111000000000",
		"00000001000011110010000011110001000011110000000111110000000011110001000000010000000100010000000000000000000000010010000000000010000000000000000100000001000000000000000011110000111100000000000100000000000000100000000100001111001000000000000100000001000000000001000000011110000100000001111100000001111100000000000000001110000011110000000011110001111100000000000111010001000000000000001100000000111100001111000000000000000000010000000000000000000000001111000100000000000011110001000011110000111111100000000000001111",
		"11110000000000000000000000000000001011111111000100000000000000000000000100000000001000000000111100010000000000000010111000000000000000000000000011110000000100010000000000000000000011110001000000010000000100010000000000001111000100010000000000000000111100000000000000001111111100011111000000110000000000000001000100000001000000000000000111110000111000000000000100000000000000000000000100000001111111110000000000000000000000001111000100000000111100001111000100001110111111101111000000001110000000000001000000010000",
		"00000000000000000001000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000010000000000000000000000001111000000000000000100000000000000000000000011110000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000100000000000011110000000000001111000000000000000011111111000000000000000100001111000000000000",
		"00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"11110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"11110001111100010000000100000000111100000001000000000000000011110001111100010000000000010000001000000001000000101111000000000001000000100000000100000000111100000000000011110000000011111111000111100001000000001111000000000010111100000001000000010001000000000000000000000000000000000000000000000001000000010000000100000001000000000000111100000000000000000000000011111111000011110000000011110000000000000000111111110000000000001111000000000000000100000001000000000000000000000000110100000000000000000000110100000000",
		"11110001000000010000000100000010111100000001000000000000000100000001000000000000111100001111001000000001111100011110000000000010000100100000000000000001111100000000000011100000000011101111000011110001111111111111000000000010111100000001000000000001000011110001111100001111000011110000000000000001000000010000000000000001000000000001111011110000000011110000000111101111000011101111000000000000000000000000111111111111000000001111000100001111001000000001000000000001000100000000110100000001000111111111111000000000",
		"00000000000100100000000100000000000111110001000000001111000100010000000000000001000000010000000000000001000000000000111111110010000000000001000000000001000000000000000100010000000011110001000000000001111000000000000000010000000000010000000000000001000011110000111100000000000000000000000000000000000000011111000000000000000100100000000011100000000011111111000011100000000011110000000000000000000000000000000000010000000011110000000100001111000111110001000000010001000100000001111111100001000011111111000011110000",
		"00000000000100010000000100000000000011110010000000000000000100000000000000010000111100011111000000000001111100000000000000000001001000000001111100000001000000000010000100000000000011110000000000000001111111100000111100000000000000100001000000100001000011110000111000001110000011110000000000000000000000010000000000010001000100010001111100000000000000001110000011111111000011100000111100000000111100000000111100000000001011111111000000000000000100000000000000010000000000000001111111110001000011110000000000000000",
		"11100000000100000000000000000000000000000011111100000000000100000001000000000000000000000000000000000000000011110001000000000001000100000001111000000010111100000010000100001110000011110000111100000000111100000011000000000000111100010001000100000001000100000000000000000000000000000010000000000000000000000000000000100001000000000010000000000001000000001111000011111110000011100001111100000000111100000001111100000000001011111110000100000000000100000001000100000000000000010000111000000001111011111110000100000001",
		"11010001000000010000000000000000000000100010000000010000000100000001000000000000000000010000111100000000000000000001000000000001000000000000000000000010000000000001000000001111000000000000111000000000110100000100000000000000111100010000000000010000000000000000111000000000000000000001000000000000111100000000000000100000000000010010000000000001000000000000000011111111111111110000000000000000000000000001000000000000000100000000000100000000000111110000000100000000000000010000000000000000111100000000000100000001",
		"11110001000000000000000000000001000011110010111100000000000000010000000000010001000000000000111111110000000000000001000000000001000000000000111100000001000000000001000000000000000100000000110100000001111011110010000100000000000000000000000000010001000000000000111100001111000000000000000000000000000000001111000000100000000000000000111100000001000000001111000000000000000100000000000100000000000000000000111100010001000000000001111100010000000100000000000100000000001000010001111100000000000000000000000100010000",
		"00000010000000000000000100000001000000000010111100000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000001111100010000000000001111001000000000000000000001110111110001000100010000000000000000000000010001000000000000111100001111000000000000000000000000000000000000000000100000000000000000000000000001000000001111111100000000000000000000000100000000000100000000000000000001000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000010000",
		"00000000000100000000000100001111000000000000111100000000000000010000000000000000111100000000000000000000000011110000111100010001000100000000111100000011000000000000000100001101000011110000111011110000110100010001000000010000000000000010000000000000111100000000110000000000111100000001000000010000000000000000111100010000000000010001000000000000000000001111000100000000000000000000000011110001111100000000000000010001000111111111000000001111000000000010000000001111000000010000111111111111111100000000000000000001",
		"00000011000000000000000000001111000100001111000000000000111100010000000100100000000000000000000000000001000111110000111100000001000011111111111100000011000000000000000100001110000000000000111100000000111100010001000000010000000000010000000000010000000000000000110100000000000000000000000000000000111100001111000000000000111100000000000000000001000000000000000011110001000000010000000100000000000000010000000000100000000011100000000100001111000000000001000011111111000100000000000000000000111000000000000000000001",
		"00000010000000000000000000000000000100000000000000000000000000000000000100100000000000000000000011110000000000000000000011110000000000001111111100000001000000000000000000001110000000000000000000000000000100010000000000010000111100010000000100010000000000000001111000000000000000000000000000000000111100000000000000000000111100000000000000000001000000000000000000000001000000000000000011111111000000010000000000100000000011110000000000000000000000000000000000001111000000000001111100000000111111110000000000000001",
		"00010010000000000000000100000000000100000000000100000000000000000001000000010001000000000000111100000000111011110000000011100001000000001111111100000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000110000111100000000000011110000000000000000000000001111000011111111000000000000111000000000000000010001000000010000000011110010000000010000000000000000000000001111000000100001000011101111000100000000000000000001000000001111000000000010000000000000000000000000111100000001",
		"00010011111111110000000100000000000111110000000000000001111100000010000000100000000000000001000000000000111000000000111000000000000000011111111000000001000000010000000000001111000011110000000000000000111100000000000000000000111100000000000000010000111000000000000011110000000000000000111100000000000100000000000000000000110100000000000100010001111100010001000011110001000000010000000000000001000000000000111100010000000011111100000000000000000000000010000000000000000000000010000000001111000000000000000000000000",
		"00000001000000000000000000000000000111110000000000000000110100000000000100110001111100010000111100000001111111110001000011110000000100011111111100000001000000000000000100001111000011110000000000000000000000000000000000000000000000010000000000010000111100000000111011110000000000000000111100001111000100000000000100000000111100000000000000000000111100010001000011110001000000000000000100000000000000000000111100010000000011111111000000000000000000010001000000000000000000000001000000000000000000001111000000010000",
		"00010011000000000000111111100000000000000000000000000000111000000000000000110000000000010001000000010001111111100001111100000000000100011111111100000000000000000000000000001111000000000000000100001111000000010000000011110000111100010000000000100000111011110000111011110000000000000000000000000000000000000000000100001110111111110000000100001111000000000001000011110001111100000000001000000001000000001111000000000010111100000000000000000000000000000001000100000000000000010001111100000000111100001111000000000000",
		"00000011000000000000111111111110000011111111000000000000111100010001000000110000000100000000000000010010111100000001000000010001000000001111000000000000000100010000000100001110000011110001000100000000000000000001000100001111111100010000000000100000000000000000111011100000111100001111111100000001000000000000000000001110000000000000000111100000111100000000000011110010000000001110000000000000111100000000000000000000111100001111000000000000000100000001000111110000000000010001000000000000111000000000000000000000",
		"00000001000100010000000000000000000000000000111100000000111100000010000000010000000000000000000000000000111100010010111000000001000000010000000000000000000000000001000000001110000000000001000100000000000000000001000000001111111100000000000100010000000000000000111100000000000000000000111100010000000100000000111100001111111100000000000011100000111111110001000000000000000000001111001000000001111100000000000100000000000000001111000100000000000011110000000011100000000000000001111100000000111100000000000000000000",
		"00000001000000000000000011110000000000000001000000000000111100000001111100010000000000010010000000010001111100000010111000000000000000010000001011110000111100010001111100001110000000000000000000000000000011110001000000001111111100000000000100000000111100000000000000001111000100000000000000100000000011110000111000000000111111110000000000000000111100000000000011100000000000001111001011110000000000011111000100000000111100000000000000000000000000000000000000001111111100000000000000000000111111110000111100000000",
		"00010000000000000000000011100000000000000000000000000000111111110000000000010000000000010000000000110000000000000001111100000001000000100000000100000000000000000001111011110000000000000010000011110000000011110001000000001111000000001111000100000000111100000000000000001111000100000000000100101111000000000000000000001111111100000000000011110000000000010000000011010000111100001111000100000000000000000000000100001111111100000000000000010000000000000000000011110000000000000000000011110000000011100000110100010000",
		"00000000000000000000111111110000000000000000000100001111000000000001000000000001000000001111000000010000000100010000000000000001111100100000000000000000000000000000111111110000000000000000000000000000000000010000000000000000000100000000000100000000000011110001000000000000000000000000000100010000000000000000000000000000111100001111000111110000000000000000000011100001000000001111000100000000000000000000000100000000111100000001000000000000111100001111000011100000000111110001000011110000000011110000111100010000",
		"11110000000000001111000011110000000000000000000100010000000000000000000000000000000100000000000000010000000100000001000000000001000000000000000000000000000000010000000011110000000000000001000000000000000000000001000000001111000100000000000000000000000000000000000000001111000000000000000000011111000000000000000000000000000000000000001011110000111100000000000011110000000000001111000000000000000000000000000000000000111100000000000000000000000000001111000011111111000000000000000011111111000011110001000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000111000000000000011110010000000010000000100000000000000010000000000000000000000001111000100000000000000100000111100100000000011110000000000010000000011110000000000000001000100000000001000000000000000001110000000000001000000000000000000000000000111110001000000011111000011110000000000000000000000000000000000010000000011110000000000010000000100000000000011110000000000001111000000001110000000001111000000001111111100011111111100000001000000001111111000000010000100000000000011110000000111100000000000000000",
		"00000000111100000000000011100011000000000000000111111111000100010000000000000001000000011111001000000001000000001111000000010010000000000001000000010010000011110000000000000001000000000000001000000001000000001110000000000001111111110000000000000001001011110010000000101111000111110000000000000000000000000001000000010000000000000000000011110001000100000001000111100000000011111111000000001110000000001111000000001110111000000000111111110000000100000000111000000010000011110000000011100000000111100000000111110000",
		"00000000000000000000000011100010000000000001000011111111000000000000000000000001000000010000001000000010000000000000000000000001000000000000000000000001111011110000000011110000000011110000000100000001111100001111000000000010000011110000000000000001000111110010000000111110000011100000000000000000000000000000000000010001000000000001000011110001000100000000000011100000111111111111000100001111000011111111000000001110111100010000000011110000001000000000111100000010000011110000111111100000000111101111000011110001",
		"11110001000000000001000100000001000000000010000011100000000000000000000000000000000000001111000000000000111000000000000000000000000100000000000000000010111100000000000000001111000011101111000000010001000000000000000000000001000011110001000100000010000000000010111100101111111100000001111100000001000111110001111100000010111100000010000100010001000000000000000111100000000011110000000100000000111011100000000000000000000000001111000011110000000100000000000000000000000000000000000000000000000011101111000011110000",
		"00000000000000000000001000000001000000000010000000000010000000000000000000000000000100000000000000010000111100000000000000000000000000000000000000000001111100000001000000001111000011110000000000010001111100000000000000010000000111110001000000000010000000000000000000000000000000100000111100010000000011110000111100000000111000000001000100000001000100000001000000001111000000000000001000000000000011110000000011110000111100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001",
		"11110001111100000000000100000001000000000001000000000010000100000000111100000000000000001111000000010000111100001111000000000000000100001111000000000001111000000001000000001111000011100000111100010001111011110001000000010000111100000000000000000011111100100001111100000000000000100001111100010000000111100001000000000000111000000001000000000001000000000000000000011111111111110000001100000000000000001111000011101111000000000000000000000000000100000000111100010000000111111111000000000000111000000000000100000001",
		"11110000000000000000000000000000000000000000111100000010000000000000000000000000000000001111000000000000000000000001000000000001000000000000111100000010000000000000000111101111000011100000111000010010111000000001000100010000000000000000111100000011000000100000111100000000000000110000000000000000001000000000000000010000111100000000111111100000000011110000000000100000000011111111000100010000000011110000111111110000000100000000000011110000000000010000111100000000000000000000111111110000111000000000000000000001",
		"00000001000000000001000000000000000011110001111100000001111100010000000000000000000100001111000000000000000000000001000011100010000000000000111100000000000000000000000111111111000000000000000100000001111000000000000100000000000100000000000000000001000000010000000000001110000000000000000000000000000100000000000000000000111100000000000011100000111111110000000000000000111100000000000000000000111100000000111100000000111100000000000000000010000000000000000000000000000000000000000011110000000000001111111111110001",
		"00000010000011110000000111110000000111100010111100000001000000000000000000100000001000010000000000000001111111100000000000000001000000001111111100000001000000010000000011110000000011110000000100000000000011110000000000000000000100000000000000000001000000100000111100000000000000000000111100010000001000000000000000010000111011110000000100000001111011100000000011110000111100001111001000000000111000000000111100000000000000001111000000000000000000000000111100010000000000000000000100000001111111110000000000000001",
		"00000010000000000000000000000000000011100000000000010010000000000001000000010000000100000000000000010001111011110000000000000001000000010000000000000000000000100001000011110000111111110000000000010001111011110010000000010000111100010000000000010001111000100000111100001110000000000000111100010000000100000000000000010000111011110001000011110000111011110000000000000001111100000000000100000000111000000000000000000000000011111110000100000000000000010001000000011111000000001111000000000000111111110000000000010010",
		"11110011000000000000000000000010000011110000000100000010000000000001111000010000000000000000000000100001111100000001000011110001000000100000111000000001111000000000000111101110111111100000111100010001111111100001000100010000000000000000000000010011111000100001111100011110000000000001000000000000000000000000000100010000111011110010000011110001110100000000000011110001111100000000001000000000111000001111111100000001000000001101000011110000000000000000000000000000000000001111111100000000111111110000000000000011",
		"11110001000000000000000000010001000000001111001000010010000000000000111100000000000000010010000000100001111100000000000011110000000000011111111000000001000000000000000111101101111100000000111100000000111111110000000100000001000000010000000000010000111000010000111100000000000000000000000000000000000000000000000100011111111100000000000111110001111100000001000011110001111000000000001000000000111111110000000000010001000011101111000000000000000000000001000000000000000000000000111000000000111000000000111100000010",
		"00000001000000000000000000000000000100000001000100000001000000000010111100000000000000000001000000010000111000000000000000000001000000111111000000000010000000010000000011111110111111110000000000010000111000000000000100010000000000000000000000000000111100010000111000000000000000000000111100000000000000000000000000011111111100000000000011110001111000000010000011110000111100001111001000000000000000000000111100000001000000001110000000000000000100000001000000000000000000010000000000000000111111110000111111110010",
		"00000001000000000000000000000000001000000010000000000010000000000001000000000000000000000000000000000001111100000000111111100001000100011111000000000001000000000000000000000000111111100001000000010001000000000000000000010000000011110000000000000001111100100000111100001110000000000001111111110000000000000000000000101111111100000000000111110001111000000001000100000000111100001111001011100000111100000000111100000001000011111111111100000001000100010000000000011111000000100000000000000000111100000000000000000001",
		"00000000000000010000000000000000000000000010000000000000000000000000000000000000000000010001000000000000111000000000111100000000000100010000111100000000000000000000000000001111000000000000111100000000001000000001000000000000000000000000111100000000000000010000111100001110000000010000111100000000000000000000000000101110111100000000000111110000111100000001000000000000000000001111000000000000111100000000000000000001000000001111000000000000000000010000000000001111000000010000000000000001111100000000000000000001",
		"11110001000100000000000100000000000000000001000000000000000000000000000000101111000000010001000000010001111100001110000000000001000100000000000000000001000000100001000100001111111011110000111100000000000000000001000100100000111100010001000000000000000000100000000000001111111100010010111000010000001000000000000000011111111100000000000011111111111100000000000000000000000000000000000000000001111100000000000000000000111000001110000011100000000000010001000000001111000000001111000000010000111000000001000000010001",
		"11110001000100000000000111110000000011110001000000000000000000000000111100100000000000000000000000100001111100010000000000000010000100010000000011110001111100010000000011111110111011110000000000010001000011110001000100010000000000000000000011110001000000110000000000001110111100000001111000000010000100000001000000101111000000000001000011110000110100000000000100000000111100001111000000000001111000001111000011110000111100011111000000000000000000000001111100001111000000000000111100000000111111110000000000010001",
		"00000000000000000000000100000000000011110001111100000000000011110000111000100000000000000001000000100001111100010000111100000001000100011111000000000001111100010000000000001110111011110000111100010000000000000001000100000000000000000000000000000001111100010000000000001110000000000010111100010001000000000001000000010000111111110001111100000000111000000000000011110000111100001111000100000000111000001111000011110000111000000000000000000000000100000000000000011111000000001111111100000000111111110000000000000001",
		"00000000000100000000000000000000000000000000000000000000000000000000000000010000000000010001000000010001000000000000000000000000000100001111000000000001000000000001000000001111111111110000000000010000000000000000000000000000111100000000000000000000111100010000000000001111000000000001111100010000000000000001000000000000000011110000111100000000111100000000000000000000000000000000000100001111000000000000000011110000111100001111111100000000000000000000000000011111000000000000000000010000111111110000000000000001",
		"00000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000100000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000001000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000111100000000000000000000111100000000111100000000000000000000000100000000000000000000000000000000000000000000000000001111000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000111100000000111100001111000011110000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000111100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00011111000100001110000000000000000011110000000000001111000011110000111100001110111100000010000000010000000000001111000100001111000100011111000100000000000000000000000000000000111100001111000011110000111100000001000000000000000000000001000000000000111100000000000011111111000000000001000000011110000100000000111111110001111000010000000000011111000100000000000000100000000100000001000000010001000100000000000011110000000100000001000000000000000000000001000100001110111111110000111100010000111100000000000000000000",
		"00101110001000001101000100011110000011010001000000001110001011100001111000001101111000000011000100010001000000001110000111111101000000101110010011100000111100100001000000001111111011111101111011010010110100000010000000000010111000000001000000000000111100001111111111101101111000010010000100111110001100000011110111010010111000111111111100111111001000100000111000101110001011110011000000110010001000010001000011010001001011100011001011101111000100010011000100111101111011110000111100100000110100100000000000000001",
		"00000000000000000000000000000000111111010000000000000000000011100000111000000000000100000001000000000001000000010000000000000001000100000000000011110001111100010000000011110000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001111000000000000000000000000100000001111100000000000100000000000000000000000100000001000000000000000000000010000000000000000000000001000000000000000000010001000000000000000000000000000011110000000000000000",
		"00000000000000000000000000000000000011110000000000000000000011110000000000000000000100000000000000000001000000010000000000000000000100000000000000000001000000010000000011110000111100000000000000000001000000000001000000000000000100000000000000000000000000000000111100010000000000000000000000010001000000000000000000000000000000000000000000000000111100000000000000000000000000000000000111110000000000000000000000000000000000010000000000000000000000000000000000000000000000001111000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000111100000000000000000001000000000000000000000000000000000000000000000000000000000000111100011111000000000000000000000000000000000000000000000000000000000001000011110000000000000000000100000000000000000000000011110000000000000000000000000000000000000000000011110000000100000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000111100000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
		"00000000000100000000000000011111000000000000000000000000000111100000111100011111000000000001000000010001111111110000000000000000000000010000000000000001000000010000000000000000111111100000000000000010111111110001000000000000000000000001000000000001000000010000000011111111111100000010111100010000000111110001111100000000000000010000000000000000111100000000000000010000111100000000000000000000000000000000000011110000000000000000001011110000000000000001000000011111000011111110000000010000111100010010000100000000",
		"00000000000000000000000000010000000011110000000000000001000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000001000000000000000000000000000011100000000100000001111011110001000000000000000000000000000000000000000000010001111100000000000000000000111100000001000000000001111111110001111000010000000000000000111100000001000000000000111100000000000111110000000000000000000011110000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000100000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111100000000000000000000000000000000111100000001000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000001000000000000111100001111000000000000000000000000000000000000111100000000111100000000000000000000000000000000000000000000111100000000000000000000000000000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000001000000000000000000000000111100000000000000000000000011110000000000001111000000000001000000010000000000000000000000000000000000000000000000000000000000010000000000000000000011111111000000000000000011110000000000000000000000000000000000000000000000010000000000001111000000000000000000000000000000000001000000000000000000000000000000000000111100000000000000000000111100000000000000000001111100000000000011110000000000000000000100000000000000000000000000000000000000000000000000000000111111110000000000000000",
		"00000001000000000000000000000000000011110000111100000001000000000001111100000000000000001111000000010000111100000000000000000001000000000000111100000000111100000000000000000000111111111111111100010001000011110000000000000000000000000000000000000000000000010000000000001110000000010001111100000000000100000001000011010000000000000001000100000000111100000000000011111111000011110000000000000000111111111111111111110000000000000000000011110000000100000000000000010000000000001111000000010000000000000000000011110000",
		"00000000111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000001000000000000000000000000000011110000000000010001001000000000000100000000000000000000000000000001000000000001111100000000000000000000000000001111000000000001111100000000111100000000000111110000111100000000000000000000111100000000000100000000000011110000111100000000000011110000000000000000000000000000000000000000000000010000000000000001000000001111000000000000",
		"00000000000000001111000000000000000000000000000000000000000011110000000000000000000000000000000000010000000000001111000000000000000000010000000000000000000000010000000000000000111111100000111100000000000000000000000000000000111100000001000000000000000000000000000000000000000000000001000000001111000000000000111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000010000000000001111000000000000000000000000111100010000000000000000",
		"00000000000100000000000000000000111100000000111100000000000011100000000000000000000000000000000000000001000000000000000000000000000000000000111100000000000000000000000000000000111111101111000000000000000000000000000000000000111100000000000000000001000000010000000000001110000000000001000000000000000100000001111000000000000000000000111100000000111100010000000000000000111100000000000000000000000000001111000011110000000000001111000000000000000100010000000000000000000000000000000000010001000000000000000000000000",
		"00000001000000000000000000000000000000000000000000000000111100000001111100000000000000000000000000000000111100000000000000000000000000000000111000000000000000000000000000000000111111101111000000010000000011110000000000000000000000000000000000000001000000010000000000001110000000010001000000000000000100000000000000000000000000000001000000000000111100000000000011110000111011110000000000000001000000000000000011110000000000001111000011110000000100000000000000000000000000001111000000010001000011110000000100000000",
		"00000000000100000000000000000001000000010000000000000000000000000000111100000000000000000000000000010000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000011110000000100000000000000000000000000000000000000001111000000000000000000000000000000010000000000000000000000000000000000000000000100000000",
		"00000000000100000000000000000000000000000001000000000000000000000000111100000000000000000000000000010000000000001111000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011110000000000000000000000000000000000000000000011110000000000001111000000001111000000000000000000000000000011110000000000000000000000000000000000000000000000000001000000000000000000000000",
		"00000000000100000000000100000000000000000001111100000000000011110001111100010000111100000000000000000001000000001111000000001111000100001111000000000000111100010001000000001111111100001111111100010000000000000000000100000000111100000000000000000001000000001111000000000000000000000001000000000000000000000001000000000000000011100000000000000000111100000000000000000000000011110000000000010000000000001111000011110000000000000001000011110000000100000000000000011111000000000000111100000001000000000000000000000000",
		"00000000000100000000000011111111000000000001000000000000000000000000000000000000111100000010000000010010000000000000000000001111000100001111000000000001111100010001000000001111111111111111000000010001000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000001000000000000000011100000000000000000000000000000000000000000000000000000000000001111000000000000000011110000111100000000111111110000000000000000000000011111000000010000000000010000000011110000000000000000",
		"00000000000100000000000000000000000011110001000000010000000000000000000000000000111100000000000000000000000000000000000000000000000000001111000000000000111100000000000000001111000000000000111100000000111100000000111100000001000000000000000000000000111100000000000000000000000000000000000000000000000100000000000000000000000000011111000000000000000000000000111100000000000011110000000100000000000100000000000011110000000011110000000000000000000100000000000000001111111100000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
	);

begin

	rom_behavior	: process(clka)
	begin

		if clka'event and clka = '1'
		then

			douta <= mem(to_integer(unsigned(addra)));

		end if;

	end process rom_behavior;

end architecture behavior;
